fp2int_inst : fp2int PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
