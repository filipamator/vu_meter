sqrt_inst : sqrt PORT MAP (
		radical	 => radical_sig,
		q	 => q_sig,
		remainder	 => remainder_sig
	);
