library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity hannwindow is
port (
        i_sample    : in STD_LOGIC_VECTOR(9 downto 0);
        o_value     : out STD_LOGIC_VECTOR(31 downto 0)
);
end hannwindow;



architecture Behavioral of hannwindow is

signal r_sample : integer range 0 to 1023 := 0;


begin


r_sample <= to_integer(unsigned(i_sample));

with r_sample select o_value  <=
    "00000000000000000000000000000000" when 0,      -- 0.0
    "00110111000111100011100011011000" when 1,      -- 9.430769E-6
    "00111000000111100011100001110111" when 2,      -- 3.7722722E-5
    "00111000101100011111111011001110" when 3,      -- 8.487479E-5
    "00111001000111100011011011101111" when 4,      -- 1.5088519E-4
    "00111001011101110011010000001100" when 5,
    "00111001101100011111101011110000" when 6,
    "00111001111100100011110110101111" when 7,
    "00111010000111100011000011010011" when 8,
    "00111010010010000011001100001110" when 9,
    "00111010011101110010010100100000" when 10,
    "00111010100101011000001101001011" when 11,
    "00111010101100011110101101111000" when 12,
    "00111010110100001100101011010001" when 13,
    "00111010111100100010000100001000" when 14,
    "00111011000010101111011011100110" when 15,
    "00111011000111100001100001100011" when 16,
    "00111011001100100111010011001010" when 17,
    "00111011010010000000101111101010" when 18,
    "00111011010111101101110110001101" when 19,
    "00111011011101101110100101111010" when 20,
    "00111011100010000001011110111011" when 21,
    "00111011100101010101011110100010" when 22,
    "00111011101000110011010001010001" when 23,
    "00111011101100011010110110100101" when 24,
    "00111011110000001100001101111010" when 25,
    "00111011110100000111010110101100" when 26,
    "00111011111000001100010000010011" when 27,
    "00111011111100011010111010000111" when 28,
    "00111100000000011001101001101111" when 29,
    "00111100000010101010101101110111" when 30,
    "00111100000101000000101001000101" when 31,
    "00111100000111011011011011000001" when 32,
    "00111100001001111011000011010011" when 33,
    "00111100001100011111100001100011" when 34,
    "00111100001111001000110101011000" when 35,
    "00111100010001110110111110010111" when 36,
    "00111100010100101001111100000101" when 37,
    "00111100010111100001101110001000" when 38,
    "00111100011010011110010100000001" when 39,
    "00111100011101011111101101010101" when 40,
    "00111100100000010010111100110010" when 41,
    "00111100100001111000011100001001" when 42,
    "00111100100011100000010100011111" when 43,
    "00111100100101001010100101100100" when 44,
    "00111100100110110111001111001000" when 45,
    "00111100101000100110010000111001" when 46,
    "00111100101010010111101010101000" when 47,
    "00111100101100001011011100000001" when 48,
    "00111100101110000001100100110100" when 49,
    "00111100101111111010000100101110" when 50,
    "00111100110001110100111011011101" when 51,
    "00111100110011110010001000101101" when 52,
    "00111100110101110001101100001011" when 53,
    "00111100110111110011100101100011" when 54,
    "00111100111001110111110100100010" when 55,
    "00111100111011111110011000110011" when 56,
    "00111100111110000111010010000001" when 57,
    "00111101000000001001001111111011" when 58,
    "00111101000001010000000001000000" when 59,
    "00111101000010010111111100000010" when 60,
    "00111101000011100001000000111000" when 61,
    "00111101000100101011001111010101" when 62,
    "00111101000101110110100111001111" when 63,
    "00111101000111000011001000011010" when 64,
    "00111101001000010000110010101010" when 65,
    "00111101001001011111100101110010" when 66,
    "00111101001010101111100001101000" when 67,
    "00111101001100000000100101111110" when 68,
    "00111101001101010010110010101000" when 69,
    "00111101001110100110000111011000" when 70,
    "00111101001111111010100100000100" when 71,
    "00111101010001010000001000011100" when 72,
    "00111101010010100110110100010101" when 73,
    "00111101010011111110100111100000" when 74,
    "00111101010101010111100001110001" when 75,
    "00111101010110110001100010111001" when 76,
    "00111101011000001100101010101010" when 77,
    "00111101011001101000111000110110" when 78,
    "00111101011011000110001101010000" when 79,
    "00111101011100100100100111101000" when 80,
    "00111101011110000100000111110001" when 81,
    "00111101011111100100101101011011" when 82,
    "00111101100000100011001100001100" when 83,
    "00111101100001010100100100001011" when 84,
    "00111101100010000110011110100101" when 85,
    "00111101100010111000111011010010" when 86,
    "00111101100011101011111010001000" when 87,
    "00111101100100011111011011000010" when 88,
    "00111101100101010011011101110110" when 89,
    "00111101100110001000000010011101" when 90,
    "00111101100110111101001000101110" when 91,
    "00111101100111110010110000100001" when 92,
    "00111101101000101000111001101111" when 93,
    "00111101101001011111100100001110" when 94,
    "00111101101010010110101111110111" when 95,
    "00111101101011001110011100100000" when 96,
    "00111101101100000110101010000010" when 97,
    "00111101101100111111011000010010" when 98,
    "00111101101101111000100111001010" when 99,
    "00111101101110110010010110011111" when 100,
    "00111101101111101100100110001001" when 101,
    "00111101110000100111010101111111" when 102,
    "00111101110001100010100101111000" when 103,
    "00111101110010011110010101101011" when 104,
    "00111101110011011010100101001101" when 105,
    "00111101110100010111010100010111" when 106,
    "00111101110101010100100010111111" when 107,
    "00111101110110010010010000111011" when 108,
    "00111101110111010000011110000010" when 109,
    "00111101111000001111001010001010" when 110,
    "00111101111001001110010101001001" when 111,
    "00111101111010001101111110110110" when 112,
    "00111101111011001110000111000111" when 113,
    "00111101111100001110101101110001" when 114,
    "00111101111101001111110010101100" when 115,
    "00111101111110010001010101101101" when 116,
    "00111101111111010011010110101001" when 117,
    "00111110000000001010111010101011" when 118,
    "00111110000000101100011000110110" when 119,
    "00111110000001001110000101101111" when 120,
    "00111110000001110000000001010001" when 121,
    "00111110000010010010001011011000" when 122,
    "00111110000010110100100011111101" when 123,
    "00111110000011010111001010111011" when 124,
    "00111110000011111010000000001110" when 125,
    "00111110000100011101000011101111" when 126,
    "00111110000101000000010101011010" when 127,
    "00111110000101100011110101001000" when 128,
    "00111110000110000111100010110101" when 129,
    "00111110000110101011011110011011" when 130,
    "00111110000111001111100111110100" when 131,
    "00111110000111110011111110111010" when 132,
    "00111110001000011000100011101001" when 133,
    "00111110001000111101010101111010" when 134,
    "00111110001001100010010101101000" when 135,
    "00111110001010000111100010101101" when 136,
    "00111110001010101100111101000011" when 137,
    "00111110001011010010100100100101" when 138,
    "00111110001011111000011001001100" when 139,
    "00111110001100011110011010110011" when 140,
    "00111110001101000100101001010100" when 141,
    "00111110001101101011000100101010" when 142,
    "00111110001110010001101100101101" when 143,
    "00111110001110111000100001011000" when 144,
    "00111110001111011111100010100110" when 145,
    "00111110010000000110110000010000" when 146,
    "00111110010000101110001010010000" when 147,
    "00111110010001010101110000011111" when 148,
    "00111110010001111101100010111001" when 149,
    "00111110010010100101100001010110" when 150,
    "00111110010011001101101011110001" when 151,
    "00111110010011110110000010000100" when 152,
    "00111110010100011110100100000111" when 153,
    "00111110010101000111010001110101" when 154,
    "00111110010101110000001011001000" when 155,
    "00111110010110011001001111111001" when 156,
    "00111110010111000010100000000010" when 157,
    "00111110010111101011111011011100" when 158,
    "00111110011000010101100010000001" when 159,
    "00111110011000111111010011101011" when 160,
    "00111110011001101001010000010100" when 161,
    "00111110011010010011010111110100" when 162,
    "00111110011010111101101010000101" when 163,
    "00111110011011101000000111000001" when 164,
    "00111110011100010010101110100001" when 165,
    "00111110011100111101100000011111" when 166,
    "00111110011101101000011100110011" when 167,
    "00111110011110010011100011011000" when 168,
    "00111110011110111110110100000111" when 169,
    "00111110011111101010001110111000" when 170,
    "00111110100000001010111001110011" when 171,
    "00111110100000100000110001000101" when 172,
    "00111110100000110110101101001110" when 173,
    "00111110100001001100101110001011" when 174,
    "00111110100001100010110011111000" when 175,
    "00111110100001111000111110010011" when 176,
    "00111110100010001111001101011000" when 177,
    "00111110100010100101100001000010" when 178,
    "00111110100010111011111001010000" when 179,
    "00111110100011010010010101111101" when 180,
    "00111110100011101000110111000110" when 181,
    "00111110100011111111011100101000" when 182,
    "00111110100100010110000110011110" when 183,
    "00111110100100101100110100100110" when 184,
    "00111110100101000011100110111100" when 185,
    "00111110100101011010011101011101" when 186,
    "00111110100101110001011000000100" when 187,
    "00111110100110001000010110101111" when 188,
    "00111110100110011111011001011001" when 189,
    "00111110100110110110100000000000" when 190,
    "00111110100111001101101010011111" when 191,
    "00111110100111100100111000110100" when 192,
    "00111110100111111100001010111010" when 193,
    "00111110101000010011100000101110" when 194,
    "00111110101000101010111010001100" when 195,
    "00111110101001000010010111010001" when 196,
    "00111110101001011001110111111001" when 197,
    "00111110101001110001011100000001" when 198,
    "00111110101010001001000011100100" when 199,
    "00111110101010100000101110100000" when 200,
    "00111110101010111000011100110000" when 201,
    "00111110101011010000001110010000" when 202,
    "00111110101011101000000010111110" when 203,
    "00111110101011111111111010110110" when 204,
    "00111110101100010111110101110011" when 205,
    "00111110101100101111110011110010" when 206,
    "00111110101101000111110100110000" when 207,
    "00111110101101011111111000101001" when 208,
    "00111110101101110111111111011000" when 209,
    "00111110101110010000001000111011" when 210,
    "00111110101110101000010101001101" when 211,
    "00111110101111000000100100001011" when 212,
    "00111110101111011000110101110001" when 213,
    "00111110101111110001001001111011" when 214,
    "00111110110000001001100000100110" when 215,
    "00111110110000100001111001101101" when 216,
    "00111110110000111010010101001101" when 217,
    "00111110110001010010110011000011" when 218,
    "00111110110001101011010011001010" when 219,
    "00111110110010000011110101011111" when 220,
    "00111110110010011100011001111101" when 221,
    "00111110110010110101000000100010" when 222,
    "00111110110011001101101001001001" when 223,
    "00111110110011100110010011101110" when 224,
    "00111110110011111111000000001110" when 225,
    "00111110110100010111101110100101" when 226,
    "00111110110100110000011110101111" when 227,
    "00111110110101001001010000101000" when 228,
    "00111110110101100010000100001100" when 229,
    "00111110110101111010111001011000" when 230,
    "00111110110110010011110000000111" when 231,
    "00111110110110101100101000010111" when 232,
    "00111110110111000101100010000010" when 233,
    "00111110110111011110011101000110" when 234,
    "00111110110111110111011001011101" when 235,
    "00111110111000010000010111000110" when 236,
    "00111110111000101001010101111010" when 237,
    "00111110111001000010010101111000" when 238,
    "00111110111001011011010110111010" when 239,
    "00111110111001110100011000111110" when 240,
    "00111110111010001101011011111110" when 241,
    "00111110111010100110011111111000" when 242,
    "00111110111010111111100100100111" when 243,
    "00111110111011011000101010001000" when 244,
    "00111110111011110001110000010110" when 245,
    "00111110111100001010110111001110" when 246,
    "00111110111100100011111110101100" when 247,
    "00111110111100111101000110101100" when 248,
    "00111110111101010110001111001010" when 249,
    "00111110111101101111011000000010" when 250,
    "00111110111110001000100001010001" when 251,
    "00111110111110100001101010110010" when 252,
    "00111110111110111010110100100010" when 253,
    "00111110111111010011111110011100" when 254,
    "00111110111111101101001000011101" when 255,
    "00111111000000000011001001010001" when 256,
    "00111111000000001111101110010010" when 257,
    "00111111000000011100010011010001" when 258,
    "00111111000000101000111000001100" when 259,
    "00111111000000110101011101000000" when 260,
    "00111111000001000010000001101101" when 261,
    "00111111000001001110100110001110" when 262,
    "00111111000001011011001010100100" when 263,
    "00111111000001100111101110101100" when 264,
    "00111111000001110100010010100100" when 265,
    "00111111000010000000110110001001" when 266,
    "00111111000010001101011001011011" when 267,
    "00111111000010011001111100010111" when 268,
    "00111111000010100110011110111011" when 269,
    "00111111000010110011000001000110" when 270,
    "00111111000010111111100010110101" when 271,
    "00111111000011001100000100000110" when 272,
    "00111111000011011000100100111000" when 273,
    "00111111000011100101000101001000" when 274,
    "00111111000011110001100100110101" when 275,
    "00111111000011111110000011111100" when 276,
    "00111111000100001010100010011100" when 277,
    "00111111000100010111000000010011" when 278,
    "00111111000100100011011101011111" when 279,
    "00111111000100101111111001111110" when 280,
    "00111111000100111100010101101110" when 281,
    "00111111000101001000110000101101" when 282,
    "00111111000101010101001010111010" when 283,
    "00111111000101100001100100010001" when 284,
    "00111111000101101101111100110010" when 285,
    "00111111000101111010010100011010" when 286,
    "00111111000110000110101011001000" when 287,
    "00111111000110010011000000111010" when 288,
    "00111111000110011111010101101101" when 289,
    "00111111000110101011101001100000" when 290,
    "00111111000110110111111100010001" when 291,
    "00111111000111000100001101111110" when 292,
    "00111111000111010000011110100110" when 293,
    "00111111000111011100101110000101" when 294,
    "00111111000111101000111100011011" when 295,
    "00111111000111110101001001100101" when 296,
    "00111111001000000001010101100010" when 297,
    "00111111001000001101100000001111" when 298,
    "00111111001000011001101001101100" when 299,
    "00111111001000100101110001110101" when 300,
    "00111111001000110001111000101001" when 301,
    "00111111001000111101111110000110" when 302,
    "00111111001001001010000010001011" when 303,
    "00111111001001010110000100110101" when 304,
    "00111111001001100010000110000011" when 305,
    "00111111001001101110000101110011" when 306,
    "00111111001001111010000100000010" when 307,
    "00111111001010000110000000101111" when 308,
    "00111111001010010001111011111001" when 309,
    "00111111001010011101110101011101" when 310,
    "00111111001010101001101101011001" when 311,
    "00111111001010110101100011101100" when 312,
    "00111111001011000001011000010100" when 313,
    "00111111001011001101001011001111" when 314,
    "00111111001011011000111100011011" when 315,
    "00111111001011100100101011110111" when 316,
    "00111111001011110000011001100000" when 317,
    "00111111001011111100000101010101" when 318,
    "00111111001100000111101111010100" when 319,
    "00111111001100010011010111011010" when 320,
    "00111111001100011110111101101000" when 321,
    "00111111001100101010100001111001" when 322,
    "00111111001100110110000100001110" when 323,
    "00111111001101000001100100100011" when 324,
    "00111111001101001101000010111000" when 325,
    "00111111001101011000011111001010" when 326,
    "00111111001101100011111001011000" when 327,
    "00111111001101101111010001100000" when 328,
    "00111111001101111010100111100000" when 329,
    "00111111001110000101111011010110" when 330,
    "00111111001110010001001101000001" when 331,
    "00111111001110011100011100011111" when 332,
    "00111111001110100111101001101101" when 333,
    "00111111001110110010110100101100" when 334,
    "00111111001110111101111101011000" when 335,
    "00111111001111001001000011110000" when 336,
    "00111111001111010100000111110010" when 337,
    "00111111001111011111001001011101" when 338,
    "00111111001111101010001000101111" when 339,
    "00111111001111110101000101100110" when 340,
    "00111111010000000000000000000000" when 341,
    "00111111010000001010110111111100" when 342,
    "00111111010000010101101101011000" when 343,
    "00111111010000100000100000010011" when 344,
    "00111111010000101011010000101010" when 345,
    "00111111010000110101111110011101" when 346,
    "00111111010001000000101001101001" when 347,
    "00111111010001001011010010001100" when 348,
    "00111111010001010101111000000110" when 349,
    "00111111010001100000011011010101" when 350,
    "00111111010001101010111011110110" when 351,
    "00111111010001110101011001101000" when 352,
    "00111111010001111111110100101011" when 353,
    "00111111010010001010001100111011" when 354,
    "00111111010010010100100010010111" when 355,
    "00111111010010011110110100111111" when 356,
    "00111111010010101001000100101111" when 357,
    "00111111010010110011010001101000" when 358,
    "00111111010010111101011011100110" when 359,
    "00111111010011000111100010101001" when 360,
    "00111111010011010001100110101111" when 361,
    "00111111010011011011100111110110" when 362,
    "00111111010011100101100101111101" when 363,
    "00111111010011101111100001000011" when 364,
    "00111111010011111001011001000101" when 365,
    "00111111010100000011001110000010" when 366,
    "00111111010100001100111111111001" when 367,
    "00111111010100010110101110101000" when 368,
    "00111111010100100000011010001111" when 369,
    "00111111010100101010000010101010" when 370,
    "00111111010100110011100111111001" when 371,
    "00111111010100111101001001111010" when 372,
    "00111111010101000110101000101100" when 373,
    "00111111010101010000000100001101" when 374,
    "00111111010101011001011100011100" when 375,
    "00111111010101100010110001011000" when 376,
    "00111111010101101100000010111111" when 377,
    "00111111010101110101010001001111" when 378,
    "00111111010101111110011100000111" when 379,
    "00111111010110000111100011100110" when 380,
    "00111111010110010000100111101010" when 381,
    "00111111010110011001101000010010" when 382,
    "00111111010110100010100101011100" when 383,
    "00111111010110101011011111001000" when 384,
    "00111111010110110100010101010011" when 385,
    "00111111010110111101000111111101" when 386,
    "00111111010111000101110111000011" when 387,
    "00111111010111001110100010100110" when 388,
    "00111111010111010111001010100010" when 389,
    "00111111010111011111101110111000" when 390,
    "00111111010111101000001111100101" when 391,
    "00111111010111110000101100101001" when 392,
    "00111111010111111001000110000001" when 393,
    "00111111011000000001011011101110" when 394,
    "00111111011000001001101101101100" when 395,
    "00111111011000010001111011111100" when 396,
    "00111111011000011010000110011100" when 397,
    "00111111011000100010001101001011" when 398,
    "00111111011000101010010000000111" when 399,
    "00111111011000110010001111001111" when 400,
    "00111111011000111010001010100010" when 401,
    "00111111011001000010000001111110" when 402,
    "00111111011001001001110101100011" when 403,
    "00111111011001010001100101010000" when 404,
    "00111111011001011001010001000010" when 405,
    "00111111011001100000111000111001" when 406,
    "00111111011001101000011100110100" when 407,
    "00111111011001101111111100110010" when 408,
    "00111111011001110111011000110001" when 409,
    "00111111011001111110110000110000" when 410,
    "00111111011010000110000100101110" when 411,
    "00111111011010001101010100101010" when 412,
    "00111111011010010100100000100011" when 413,
    "00111111011010011011101000010111" when 414,
    "00111111011010100010101100000111" when 415,
    "00111111011010101001101011101111" when 416,
    "00111111011010110000100111010001" when 417,
    "00111111011010110111011110101001" when 418,
    "00111111011010111110010001111000" when 419,
    "00111111011011000101000000111101" when 420,
    "00111111011011001011101011110101" when 421,
    "00111111011011010010010010100001" when 422,
    "00111111011011011000110100111110" when 423,
    "00111111011011011111010011001101" when 424,
    "00111111011011100101101101001100" when 425,
    "00111111011011101100000010111011" when 426,
    "00111111011011110010010100010111" when 427,
    "00111111011011111000100001100001" when 428,
    "00111111011011111110101010010111" when 429,
    "00111111011100000100101110111000" when 430,
    "00111111011100001010101111000100" when 431,
    "00111111011100010000101010111001" when 432,
    "00111111011100010110100010010111" when 433,
    "00111111011100011100010101011100" when 434,
    "00111111011100100010000100001000" when 435,
    "00111111011100100111101110011010" when 436,
    "00111111011100101101010100010001" when 437,
    "00111111011100110010110101101100" when 438,
    "00111111011100111000010010101010" when 439,
    "00111111011100111101101011001011" when 440,
    "00111111011101000010111111001101" when 441,
    "00111111011101001000001110110000" when 442,
    "00111111011101001101011001110011" when 443,
    "00111111011101010010100000010101" when 444,
    "00111111011101010111100010010101" when 445,
    "00111111011101011100011111110100" when 446,
    "00111111011101100001011000101110" when 447,
    "00111111011101100110001101000101" when 448,
    "00111111011101101010111100111000" when 449,
    "00111111011101101111101000000100" when 450,
    "00111111011101110100001110101011" when 451,
    "00111111011101111000110000101011" when 452,
    "00111111011101111101001110000011" when 453,
    "00111111011110000001100110110011" when 454,
    "00111111011110000101111010111010" when 455,
    "00111111011110001010001010011000" when 456,
    "00111111011110001110010101001011" when 457,
    "00111111011110010010011011010100" when 458,
    "00111111011110010110011100110001" when 459,
    "00111111011110011010011001100001" when 460,
    "00111111011110011110010001100101" when 461,
    "00111111011110100010000100111100" when 462,
    "00111111011110100101110011100101" when 463,
    "00111111011110101001011101011111" when 464,
    "00111111011110101101000010101010" when 465,
    "00111111011110110000100011000110" when 466,
    "00111111011110110011111110110001" when 467,
    "00111111011110110111010101101100" when 468,
    "00111111011110111010100111110110" when 469,
    "00111111011110111101110101001101" when 470,
    "00111111011111000000111101110011" when 471,
    "00111111011111000100000001100110" when 472,
    "00111111011111000111000000100101" when 473,
    "00111111011111001001111010110001" when 474,
    "00111111011111001100110000001001" when 475,
    "00111111011111001111100000101101" when 476,
    "00111111011111010010001100011011" when 477,
    "00111111011111010100110011010100" when 478,
    "00111111011111010111010101011000" when 479,
    "00111111011111011001110010100101" when 480,
    "00111111011111011100001010111011" when 481,
    "00111111011111011110011110011011" when 482,
    "00111111011111100000101101000100" when 483,
    "00111111011111100010110110110100" when 484,
    "00111111011111100100111011101101" when 485,
    "00111111011111100110111011101110" when 486,
    "00111111011111101000110110110110" when 487,
    "00111111011111101010101101000101" when 488,
    "00111111011111101100011110011011" when 489,
    "00111111011111101110001010111000" when 490,
    "00111111011111101111110010011011" when 491,
    "00111111011111110001010101000100" when 492,
    "00111111011111110010110010110011" when 493,
    "00111111011111110100001011100111" when 494,
    "00111111011111110101011111100001" when 495,
    "00111111011111110110101110100000" when 496,
    "00111111011111110111111000100100" when 497,
    "00111111011111111000111101101100" when 498,
    "00111111011111111001111101111010" when 499,
    "00111111011111111010111001001100" when 500,
    "00111111011111111011101111100010" when 501,
    "00111111011111111100100000111100" when 502,
    "00111111011111111101001101011011" when 503,
    "00111111011111111101110100111110" when 504,
    "00111111011111111110010111100100" when 505,
    "00111111011111111110110101001110" when 506,
    "00111111011111111111001101111100" when 507,
    "00111111011111111111100001101110" when 508,
    "00111111011111111111110000100011" when 509,
    "00111111011111111111111010011100" when 510,
    "00111111011111111111111111011000" when 511,
    "00111111011111111111111111011000" when 512,
    "00111111011111111111111010011100" when 513,
    "00111111011111111111110000100011" when 514,
    "00111111011111111111100001101110" when 515,
    "00111111011111111111001101111100" when 516,
    "00111111011111111110110101001110" when 517,
    "00111111011111111110010111100100" when 518,
    "00111111011111111101110100111110" when 519,
    "00111111011111111101001101011011" when 520,
    "00111111011111111100100000111100" when 521,
    "00111111011111111011101111100010" when 522,
    "00111111011111111010111001001100" when 523,
    "00111111011111111001111101111010" when 524,
    "00111111011111111000111101101100" when 525,
    "00111111011111110111111000100100" when 526,
    "00111111011111110110101110100000" when 527,
    "00111111011111110101011111100001" when 528,
    "00111111011111110100001011100111" when 529,
    "00111111011111110010110010110011" when 530,
    "00111111011111110001010101000100" when 531,
    "00111111011111101111110010011011" when 532,
    "00111111011111101110001010111000" when 533,
    "00111111011111101100011110011011" when 534,
    "00111111011111101010101101000101" when 535,
    "00111111011111101000110110110110" when 536,
    "00111111011111100110111011101110" when 537,
    "00111111011111100100111011101101" when 538,
    "00111111011111100010110110110100" when 539,
    "00111111011111100000101101000100" when 540,
    "00111111011111011110011110011011" when 541,
    "00111111011111011100001010111011" when 542,
    "00111111011111011001110010100101" when 543,
    "00111111011111010111010101011000" when 544,
    "00111111011111010100110011010100" when 545,
    "00111111011111010010001100011011" when 546,
    "00111111011111001111100000101101" when 547,
    "00111111011111001100110000001001" when 548,
    "00111111011111001001111010110001" when 549,
    "00111111011111000111000000100101" when 550,
    "00111111011111000100000001100110" when 551,
    "00111111011111000000111101110011" when 552,
    "00111111011110111101110101001101" when 553,
    "00111111011110111010100111110110" when 554,
    "00111111011110110111010101101100" when 555,
    "00111111011110110011111110110001" when 556,
    "00111111011110110000100011000110" when 557,
    "00111111011110101101000010101010" when 558,
    "00111111011110101001011101011111" when 559,
    "00111111011110100101110011100101" when 560,
    "00111111011110100010000100111100" when 561,
    "00111111011110011110010001100101" when 562,
    "00111111011110011010011001100001" when 563,
    "00111111011110010110011100110001" when 564,
    "00111111011110010010011011010100" when 565,
    "00111111011110001110010101001011" when 566,
    "00111111011110001010001010011000" when 567,
    "00111111011110000101111010111010" when 568,
    "00111111011110000001100110110011" when 569,
    "00111111011101111101001110000011" when 570,
    "00111111011101111000110000101011" when 571,
    "00111111011101110100001110101011" when 572,
    "00111111011101101111101000000100" when 573,
    "00111111011101101010111100111000" when 574,
    "00111111011101100110001101000101" when 575,
    "00111111011101100001011000101110" when 576,
    "00111111011101011100011111110100" when 577,
    "00111111011101010111100010010101" when 578,
    "00111111011101010010100000010101" when 579,
    "00111111011101001101011001110011" when 580,
    "00111111011101001000001110110000" when 581,
    "00111111011101000010111111001101" when 582,
    "00111111011100111101101011001011" when 583,
    "00111111011100111000010010101010" when 584,
    "00111111011100110010110101101100" when 585,
    "00111111011100101101010100010001" when 586,
    "00111111011100100111101110011010" when 587,
    "00111111011100100010000100001000" when 588,
    "00111111011100011100010101011100" when 589,
    "00111111011100010110100010010111" when 590,
    "00111111011100010000101010111001" when 591,
    "00111111011100001010101111000100" when 592,
    "00111111011100000100101110111000" when 593,
    "00111111011011111110101010010111" when 594,
    "00111111011011111000100001100001" when 595,
    "00111111011011110010010100010111" when 596,
    "00111111011011101100000010111011" when 597,
    "00111111011011100101101101001100" when 598,
    "00111111011011011111010011001101" when 599,
    "00111111011011011000110100111110" when 600,
    "00111111011011010010010010100001" when 601,
    "00111111011011001011101011110101" when 602,
    "00111111011011000101000000111101" when 603,
    "00111111011010111110010001111000" when 604,
    "00111111011010110111011110101001" when 605,
    "00111111011010110000100111010001" when 606,
    "00111111011010101001101011101111" when 607,
    "00111111011010100010101100000111" when 608,
    "00111111011010011011101000010111" when 609,
    "00111111011010010100100000100011" when 610,
    "00111111011010001101010100101010" when 611,
    "00111111011010000110000100101110" when 612,
    "00111111011001111110110000110000" when 613,
    "00111111011001110111011000110001" when 614,
    "00111111011001101111111100110010" when 615,
    "00111111011001101000011100110100" when 616,
    "00111111011001100000111000111001" when 617,
    "00111111011001011001010001000010" when 618,
    "00111111011001010001100101010000" when 619,
    "00111111011001001001110101100011" when 620,
    "00111111011001000010000001111110" when 621,
    "00111111011000111010001010100010" when 622,
    "00111111011000110010001111001111" when 623,
    "00111111011000101010010000000111" when 624,
    "00111111011000100010001101001011" when 625,
    "00111111011000011010000110011100" when 626,
    "00111111011000010001111011111100" when 627,
    "00111111011000001001101101101100" when 628,
    "00111111011000000001011011101110" when 629,
    "00111111010111111001000110000001" when 630,
    "00111111010111110000101100101001" when 631,
    "00111111010111101000001111100101" when 632,
    "00111111010111011111101110111000" when 633,
    "00111111010111010111001010100010" when 634,
    "00111111010111001110100010100110" when 635,
    "00111111010111000101110111000011" when 636,
    "00111111010110111101000111111101" when 637,
    "00111111010110110100010101010011" when 638,
    "00111111010110101011011111001000" when 639,
    "00111111010110100010100101011100" when 640,
    "00111111010110011001101000010010" when 641,
    "00111111010110010000100111101010" when 642,
    "00111111010110000111100011100110" when 643,
    "00111111010101111110011100000111" when 644,
    "00111111010101110101010001001111" when 645,
    "00111111010101101100000010111111" when 646,
    "00111111010101100010110001011000" when 647,
    "00111111010101011001011100011100" when 648,
    "00111111010101010000000100001101" when 649,
    "00111111010101000110101000101100" when 650,
    "00111111010100111101001001111010" when 651,
    "00111111010100110011100111111001" when 652,
    "00111111010100101010000010101010" when 653,
    "00111111010100100000011010001111" when 654,
    "00111111010100010110101110101000" when 655,
    "00111111010100001100111111111001" when 656,
    "00111111010100000011001110000010" when 657,
    "00111111010011111001011001000101" when 658,
    "00111111010011101111100001000011" when 659,
    "00111111010011100101100101111101" when 660,
    "00111111010011011011100111110110" when 661,
    "00111111010011010001100110101111" when 662,
    "00111111010011000111100010101001" when 663,
    "00111111010010111101011011100110" when 664,
    "00111111010010110011010001101000" when 665,
    "00111111010010101001000100101111" when 666,
    "00111111010010011110110100111111" when 667,
    "00111111010010010100100010010111" when 668,
    "00111111010010001010001100111011" when 669,
    "00111111010001111111110100101011" when 670,
    "00111111010001110101011001101000" when 671,
    "00111111010001101010111011110110" when 672,
    "00111111010001100000011011010101" when 673,
    "00111111010001010101111000000110" when 674,
    "00111111010001001011010010001100" when 675,
    "00111111010001000000101001101001" when 676,
    "00111111010000110101111110011101" when 677,
    "00111111010000101011010000101010" when 678,
    "00111111010000100000100000010011" when 679,
    "00111111010000010101101101011000" when 680,
    "00111111010000001010110111111100" when 681,
    "00111111010000000000000000000000" when 682,
    "00111111001111110101000101100110" when 683,
    "00111111001111101010001000101111" when 684,
    "00111111001111011111001001011101" when 685,
    "00111111001111010100000111110010" when 686,
    "00111111001111001001000011110000" when 687,
    "00111111001110111101111101011000" when 688,
    "00111111001110110010110100101100" when 689,
    "00111111001110100111101001101101" when 690,
    "00111111001110011100011100011111" when 691,
    "00111111001110010001001101000001" when 692,
    "00111111001110000101111011010110" when 693,
    "00111111001101111010100111100000" when 694,
    "00111111001101101111010001100000" when 695,
    "00111111001101100011111001011000" when 696,
    "00111111001101011000011111001010" when 697,
    "00111111001101001101000010111000" when 698,
    "00111111001101000001100100100011" when 699,
    "00111111001100110110000100001110" when 700,
    "00111111001100101010100001111001" when 701,
    "00111111001100011110111101101000" when 702,
    "00111111001100010011010111011010" when 703,
    "00111111001100000111101111010100" when 704,
    "00111111001011111100000101010101" when 705,
    "00111111001011110000011001100000" when 706,
    "00111111001011100100101011110111" when 707,
    "00111111001011011000111100011011" when 708,
    "00111111001011001101001011001111" when 709,
    "00111111001011000001011000010100" when 710,
    "00111111001010110101100011101100" when 711,
    "00111111001010101001101101011001" when 712,
    "00111111001010011101110101011101" when 713,
    "00111111001010010001111011111001" when 714,
    "00111111001010000110000000101111" when 715,
    "00111111001001111010000100000010" when 716,
    "00111111001001101110000101110011" when 717,
    "00111111001001100010000110000011" when 718,
    "00111111001001010110000100110101" when 719,
    "00111111001001001010000010001011" when 720,
    "00111111001000111101111110000110" when 721,
    "00111111001000110001111000101001" when 722,
    "00111111001000100101110001110101" when 723,
    "00111111001000011001101001101100" when 724,
    "00111111001000001101100000001111" when 725,
    "00111111001000000001010101100010" when 726,
    "00111111000111110101001001100101" when 727,
    "00111111000111101000111100011011" when 728,
    "00111111000111011100101110000101" when 729,
    "00111111000111010000011110100110" when 730,
    "00111111000111000100001101111110" when 731,
    "00111111000110110111111100010001" when 732,
    "00111111000110101011101001100000" when 733,
    "00111111000110011111010101101101" when 734,
    "00111111000110010011000000111010" when 735,
    "00111111000110000110101011001000" when 736,
    "00111111000101111010010100011010" when 737,
    "00111111000101101101111100110010" when 738,
    "00111111000101100001100100010001" when 739,
    "00111111000101010101001010111010" when 740,
    "00111111000101001000110000101101" when 741,
    "00111111000100111100010101101110" when 742,
    "00111111000100101111111001111110" when 743,
    "00111111000100100011011101011111" when 744,
    "00111111000100010111000000010011" when 745,
    "00111111000100001010100010011100" when 746,
    "00111111000011111110000011111100" when 747,
    "00111111000011110001100100110101" when 748,
    "00111111000011100101000101001000" when 749,
    "00111111000011011000100100111000" when 750,
    "00111111000011001100000100000110" when 751,
    "00111111000010111111100010110101" when 752,
    "00111111000010110011000001000110" when 753,
    "00111111000010100110011110111011" when 754,
    "00111111000010011001111100010111" when 755,
    "00111111000010001101011001011011" when 756,
    "00111111000010000000110110001001" when 757,
    "00111111000001110100010010100100" when 758,
    "00111111000001100111101110101100" when 759,
    "00111111000001011011001010100100" when 760,
    "00111111000001001110100110001110" when 761,
    "00111111000001000010000001101101" when 762,
    "00111111000000110101011101000000" when 763,
    "00111111000000101000111000001100" when 764,
    "00111111000000011100010011010001" when 765,
    "00111111000000001111101110010010" when 766,
    "00111111000000000011001001010001" when 767,
    "00111110111111101101001000011101" when 768,
    "00111110111111010011111110011100" when 769,
    "00111110111110111010110100100010" when 770,
    "00111110111110100001101010110010" when 771,
    "00111110111110001000100001010001" when 772,
    "00111110111101101111011000000010" when 773,
    "00111110111101010110001111001010" when 774,
    "00111110111100111101000110101100" when 775,
    "00111110111100100011111110101100" when 776,
    "00111110111100001010110111001110" when 777,
    "00111110111011110001110000010110" when 778,
    "00111110111011011000101010001000" when 779,
    "00111110111010111111100100100111" when 780,
    "00111110111010100110011111111000" when 781,
    "00111110111010001101011011111110" when 782,
    "00111110111001110100011000111110" when 783,
    "00111110111001011011010110111010" when 784,
    "00111110111001000010010101111000" when 785,
    "00111110111000101001010101111010" when 786,
    "00111110111000010000010111000110" when 787,
    "00111110110111110111011001011101" when 788,
    "00111110110111011110011101000110" when 789,
    "00111110110111000101100010000010" when 790,
    "00111110110110101100101000010111" when 791,
    "00111110110110010011110000000111" when 792,
    "00111110110101111010111001011000" when 793,
    "00111110110101100010000100001100" when 794,
    "00111110110101001001010000101000" when 795,
    "00111110110100110000011110101111" when 796,
    "00111110110100010111101110100101" when 797,
    "00111110110011111111000000001110" when 798,
    "00111110110011100110010011101110" when 799,
    "00111110110011001101101001001001" when 800,
    "00111110110010110101000000100010" when 801,
    "00111110110010011100011001111101" when 802,
    "00111110110010000011110101011111" when 803,
    "00111110110001101011010011001010" when 804,
    "00111110110001010010110011000011" when 805,
    "00111110110000111010010101001101" when 806,
    "00111110110000100001111001101101" when 807,
    "00111110110000001001100000100110" when 808,
    "00111110101111110001001001111011" when 809,
    "00111110101111011000110101110001" when 810,
    "00111110101111000000100100001011" when 811,
    "00111110101110101000010101001101" when 812,
    "00111110101110010000001000111011" when 813,
    "00111110101101110111111111011000" when 814,
    "00111110101101011111111000101001" when 815,
    "00111110101101000111110100110000" when 816,
    "00111110101100101111110011110010" when 817,
    "00111110101100010111110101110011" when 818,
    "00111110101011111111111010110110" when 819,
    "00111110101011101000000010111110" when 820,
    "00111110101011010000001110010000" when 821,
    "00111110101010111000011100110000" when 822,
    "00111110101010100000101110100000" when 823,
    "00111110101010001001000011100100" when 824,
    "00111110101001110001011100000001" when 825,
    "00111110101001011001110111111001" when 826,
    "00111110101001000010010111010001" when 827,
    "00111110101000101010111010001100" when 828,
    "00111110101000010011100000101110" when 829,
    "00111110100111111100001010111010" when 830,
    "00111110100111100100111000110100" when 831,
    "00111110100111001101101010011111" when 832,
    "00111110100110110110100000000000" when 833,
    "00111110100110011111011001011001" when 834,
    "00111110100110001000010110101111" when 835,
    "00111110100101110001011000000100" when 836,
    "00111110100101011010011101011101" when 837,
    "00111110100101000011100110111100" when 838,
    "00111110100100101100110100100110" when 839,
    "00111110100100010110000110011110" when 840,
    "00111110100011111111011100101000" when 841,
    "00111110100011101000110111000110" when 842,
    "00111110100011010010010101111101" when 843,
    "00111110100010111011111001010000" when 844,
    "00111110100010100101100001000010" when 845,
    "00111110100010001111001101011000" when 846,
    "00111110100001111000111110010011" when 847,
    "00111110100001100010110011111000" when 848,
    "00111110100001001100101110001011" when 849,
    "00111110100000110110101101001110" when 850,
    "00111110100000100000110001000101" when 851,
    "00111110100000001010111001110011" when 852,
    "00111110011111101010001110111000" when 853,
    "00111110011110111110110100000111" when 854,
    "00111110011110010011100011011000" when 855,
    "00111110011101101000011100110011" when 856,
    "00111110011100111101100000011111" when 857,
    "00111110011100010010101110100001" when 858,
    "00111110011011101000000111000001" when 859,
    "00111110011010111101101010000101" when 860,
    "00111110011010010011010111110100" when 861,
    "00111110011001101001010000010100" when 862,
    "00111110011000111111010011101011" when 863,
    "00111110011000010101100010000001" when 864,
    "00111110010111101011111011011100" when 865,
    "00111110010111000010100000000010" when 866,
    "00111110010110011001001111111001" when 867,
    "00111110010101110000001011001000" when 868,
    "00111110010101000111010001110101" when 869,
    "00111110010100011110100100000111" when 870,
    "00111110010011110110000010000100" when 871,
    "00111110010011001101101011110001" when 872,
    "00111110010010100101100001010110" when 873,
    "00111110010001111101100010111001" when 874,
    "00111110010001010101110000011111" when 875,
    "00111110010000101110001010010000" when 876,
    "00111110010000000110110000010000" when 877,
    "00111110001111011111100010100110" when 878,
    "00111110001110111000100001011000" when 879,
    "00111110001110010001101100101101" when 880,
    "00111110001101101011000100101010" when 881,
    "00111110001101000100101001010100" when 882,
    "00111110001100011110011010110011" when 883,
    "00111110001011111000011001001100" when 884,
    "00111110001011010010100100100101" when 885,
    "00111110001010101100111101000011" when 886,
    "00111110001010000111100010101101" when 887,
    "00111110001001100010010101101000" when 888,
    "00111110001000111101010101111010" when 889,
    "00111110001000011000100011101001" when 890,
    "00111110000111110011111110111010" when 891,
    "00111110000111001111100111110100" when 892,
    "00111110000110101011011110011011" when 893,
    "00111110000110000111100010110101" when 894,
    "00111110000101100011110101001000" when 895,
    "00111110000101000000010101011010" when 896,
    "00111110000100011101000011101111" when 897,
    "00111110000011111010000000001110" when 898,
    "00111110000011010111001010111011" when 899,
    "00111110000010110100100011111101" when 900,
    "00111110000010010010001011011000" when 901,
    "00111110000001110000000001010001" when 902,
    "00111110000001001110000101101111" when 903,
    "00111110000000101100011000110110" when 904,
    "00111110000000001010111010101011" when 905,
    "00111101111111010011010110101001" when 906,
    "00111101111110010001010101101101" when 907,
    "00111101111101001111110010101100" when 908,
    "00111101111100001110101101110001" when 909,
    "00111101111011001110000111000111" when 910,
    "00111101111010001101111110110110" when 911,
    "00111101111001001110010101001001" when 912,
    "00111101111000001111001010001010" when 913,
    "00111101110111010000011110000010" when 914,
    "00111101110110010010010000111011" when 915,
    "00111101110101010100100010111111" when 916,
    "00111101110100010111010100010111" when 917,
    "00111101110011011010100101001101" when 918,
    "00111101110010011110010101101011" when 919,
    "00111101110001100010100101111000" when 920,
    "00111101110000100111010101111111" when 921,
    "00111101101111101100100110001001" when 922,
    "00111101101110110010010110011111" when 923,
    "00111101101101111000100111001010" when 924,
    "00111101101100111111011000010010" when 925,
    "00111101101100000110101010000010" when 926,
    "00111101101011001110011100100000" when 927,
    "00111101101010010110101111110111" when 928,
    "00111101101001011111100100001110" when 929,
    "00111101101000101000111001101111" when 930,
    "00111101100111110010110000100001" when 931,
    "00111101100110111101001000101110" when 932,
    "00111101100110001000000010011101" when 933,
    "00111101100101010011011101110110" when 934,
    "00111101100100011111011011000010" when 935,
    "00111101100011101011111010001000" when 936,
    "00111101100010111000111011010010" when 937,
    "00111101100010000110011110100101" when 938,
    "00111101100001010100100100001011" when 939,
    "00111101100000100011001100001100" when 940,
    "00111101011111100100101101011011" when 941,
    "00111101011110000100000111110001" when 942,
    "00111101011100100100100111101000" when 943,
    "00111101011011000110001101010000" when 944,
    "00111101011001101000111000110110" when 945,
    "00111101011000001100101010101010" when 946,
    "00111101010110110001100010111001" when 947,
    "00111101010101010111100001110001" when 948,
    "00111101010011111110100111100000" when 949,
    "00111101010010100110110100010101" when 950,
    "00111101010001010000001000011100" when 951,
    "00111101001111111010100100000100" when 952,
    "00111101001110100110000111011000" when 953,
    "00111101001101010010110010101000" when 954,
    "00111101001100000000100101111110" when 955,
    "00111101001010101111100001101000" when 956,
    "00111101001001011111100101110010" when 957,
    "00111101001000010000110010101010" when 958,
    "00111101000111000011001000011010" when 959,
    "00111101000101110110100111001111" when 960,
    "00111101000100101011001111010101" when 961,
    "00111101000011100001000000111000" when 962,
    "00111101000010010111111100000010" when 963,
    "00111101000001010000000001000000" when 964,
    "00111101000000001001001111111011" when 965,
    "00111100111110000111010010000001" when 966,
    "00111100111011111110011000110011" when 967,
    "00111100111001110111110100100010" when 968,
    "00111100110111110011100101100011" when 969,
    "00111100110101110001101100001011" when 970,
    "00111100110011110010001000101101" when 971,
    "00111100110001110100111011011101" when 972,
    "00111100101111111010000100101110" when 973,
    "00111100101110000001100100110100" when 974,
    "00111100101100001011011100000001" when 975,
    "00111100101010010111101010101000" when 976,
    "00111100101000100110010000111001" when 977,
    "00111100100110110111001111001000" when 978,
    "00111100100101001010100101100100" when 979,
    "00111100100011100000010100011111" when 980,
    "00111100100001111000011100001001" when 981,
    "00111100100000010010111100110010" when 982,
    "00111100011101011111101101010101" when 983,
    "00111100011010011110010100000001" when 984,
    "00111100010111100001101110001000" when 985,
    "00111100010100101001111100000101" when 986,
    "00111100010001110110111110010111" when 987,
    "00111100001111001000110101011000" when 988,
    "00111100001100011111100001100011" when 989,
    "00111100001001111011000011010011" when 990,
    "00111100000111011011011011000001" when 991,
    "00111100000101000000101001000101" when 992,
    "00111100000010101010101101110111" when 993,
    "00111100000000011001101001101111" when 994,
    "00111011111100011010111010000111" when 995,
    "00111011111000001100010000010011" when 996,
    "00111011110100000111010110101100" when 997,
    "00111011110000001100001101111010" when 998,
    "00111011101100011010110110100101" when 999,
    "00111011101000110011010001010001" when 1000,
    "00111011100101010101011110100010" when 1001,
    "00111011100010000001011110111011" when 1002,
    "00111011011101101110100101111010" when 1003,
    "00111011010111101101110110001101" when 1004,
    "00111011010010000000101111101010" when 1005,
    "00111011001100100111010011001010" when 1006,
    "00111011000111100001100001100011" when 1007,
    "00111011000010101111011011100110" when 1008,
    "00111010111100100010000100001000" when 1009,
    "00111010110100001100101011010001" when 1010,
    "00111010101100011110101101111000" when 1011,
    "00111010100101011000001101001011" when 1012,
    "00111010011101110010010100100000" when 1013,
    "00111010010010000011001100001110" when 1014,
    "00111010000111100011000011010011" when 1015,
    "00111001111100100011110110101111" when 1016,
    "00111001101100011111101011110000" when 1017,
    "00111001011101110011010000001100" when 1018,
    "00111001000111100011011011101111" when 1019,
    "00111000101100011111111011001110" when 1020,
    "00111000000111100011100001110111" when 1021,
    "00110111000111100011100011011000" when 1022,
    "00000000000000000000000000000000" when 1023,       -- 0.0
    "00000000000000000000000000000000" when others;

end Behavioral;