fplog_inst : fplog PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		result	 => result_sig
	);
