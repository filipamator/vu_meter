-- megafunction wizard: %ALTFP_LOG%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_LOG 

-- ============================================================
-- File Name: fplog.vhd
-- Megafunction Name(s):
-- 			ALTFP_LOG
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 16.1.0 Build 196 10/24/2016 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2016  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Intel and sold by Intel or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--altfp_log CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" PIPELINE=21 WIDTH_EXP=8 WIDTH_MAN=23 clock data nan result zero
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" PIPELINE=1 SHIFTDIR="LEFT" WIDTH=32 WIDTHDIST=5 aclr clk_en clock data distance result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END

--synthesis_resources = reg 33 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altbarrel_shift_itd IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END fplog_altbarrel_shift_itd;

 ARCHITECTURE RTL OF fplog_altbarrel_shift_itd IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range268w280w281w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range268w276w277w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range289w301w302w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range289w297w298w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range311w323w324w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range311w319w320w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range333w345w346w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range333w341w342w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range355w367w368w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range355w363w364w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range268w272w273w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range289w293w294w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range311w315w316w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range333w337w338w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range355w359w360w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range268w280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range268w276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range289w301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range289w297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range311w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range311w319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range333w345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range333w341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range355w367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range355w363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_dir_w_range265w279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_dir_w_range287w300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_dir_w_range308w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_dir_w_range330w344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_dir_w_range352w366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range268w272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range289w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range311w315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range333w337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range355w359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range268w280w281w282w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range289w301w302w303w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range311w323w324w325w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range333w345w346w347w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range355w367w368w369w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w283w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w304w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w326w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w348w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w370w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (191 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (159 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w275w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w278w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w296w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w299w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w318w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w321w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w340w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w343w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w362w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w365w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_dir_w_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_dir_w_range287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_dir_w_range308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_dir_w_range330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_dir_w_range352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sbit_w_range328w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sbit_w_range350w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sbit_w_range263w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sbit_w_range286w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sbit_w_range306w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sel_w_range268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sel_w_range289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sel_w_range311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sel_w_range333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sel_w_range355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_smux_w_range371w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range268w280w281w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range268w280w(0) AND wire_Lshiftsmall_w278w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range268w276w277w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range268w276w(0) AND wire_Lshiftsmall_w275w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range289w301w302w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range289w301w(0) AND wire_Lshiftsmall_w299w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range289w297w298w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range289w297w(0) AND wire_Lshiftsmall_w296w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range311w323w324w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range311w323w(0) AND wire_Lshiftsmall_w321w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range311w319w320w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range311w319w(0) AND wire_Lshiftsmall_w318w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range333w345w346w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range333w345w(0) AND wire_Lshiftsmall_w343w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range333w341w342w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range333w341w(0) AND wire_Lshiftsmall_w340w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range355w367w368w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range355w367w(0) AND wire_Lshiftsmall_w365w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range355w363w364w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range355w363w(0) AND wire_Lshiftsmall_w362w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range268w272w273w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range268w272w(0) AND wire_Lshiftsmall_w_sbit_w_range263w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range289w293w294w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range289w293w(0) AND wire_Lshiftsmall_w_sbit_w_range286w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range311w315w316w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range311w315w(0) AND wire_Lshiftsmall_w_sbit_w_range306w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range333w337w338w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range333w337w(0) AND wire_Lshiftsmall_w_sbit_w_range328w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range355w359w360w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range355w359w(0) AND wire_Lshiftsmall_w_sbit_w_range350w(i);
	END GENERATE loop14;
	wire_Lshiftsmall_w_lg_w_sel_w_range268w280w(0) <= wire_Lshiftsmall_w_sel_w_range268w(0) AND wire_Lshiftsmall_w_lg_w_dir_w_range265w279w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range268w276w(0) <= wire_Lshiftsmall_w_sel_w_range268w(0) AND wire_Lshiftsmall_w_dir_w_range265w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range289w301w(0) <= wire_Lshiftsmall_w_sel_w_range289w(0) AND wire_Lshiftsmall_w_lg_w_dir_w_range287w300w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range289w297w(0) <= wire_Lshiftsmall_w_sel_w_range289w(0) AND wire_Lshiftsmall_w_dir_w_range287w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range311w323w(0) <= wire_Lshiftsmall_w_sel_w_range311w(0) AND wire_Lshiftsmall_w_lg_w_dir_w_range308w322w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range311w319w(0) <= wire_Lshiftsmall_w_sel_w_range311w(0) AND wire_Lshiftsmall_w_dir_w_range308w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range333w345w(0) <= wire_Lshiftsmall_w_sel_w_range333w(0) AND wire_Lshiftsmall_w_lg_w_dir_w_range330w344w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range333w341w(0) <= wire_Lshiftsmall_w_sel_w_range333w(0) AND wire_Lshiftsmall_w_dir_w_range330w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range355w367w(0) <= wire_Lshiftsmall_w_sel_w_range355w(0) AND wire_Lshiftsmall_w_lg_w_dir_w_range352w366w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range355w363w(0) <= wire_Lshiftsmall_w_sel_w_range355w(0) AND wire_Lshiftsmall_w_dir_w_range352w(0);
	wire_Lshiftsmall_w_lg_w_dir_w_range265w279w(0) <= NOT wire_Lshiftsmall_w_dir_w_range265w(0);
	wire_Lshiftsmall_w_lg_w_dir_w_range287w300w(0) <= NOT wire_Lshiftsmall_w_dir_w_range287w(0);
	wire_Lshiftsmall_w_lg_w_dir_w_range308w322w(0) <= NOT wire_Lshiftsmall_w_dir_w_range308w(0);
	wire_Lshiftsmall_w_lg_w_dir_w_range330w344w(0) <= NOT wire_Lshiftsmall_w_dir_w_range330w(0);
	wire_Lshiftsmall_w_lg_w_dir_w_range352w366w(0) <= NOT wire_Lshiftsmall_w_dir_w_range352w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range268w272w(0) <= NOT wire_Lshiftsmall_w_sel_w_range268w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range289w293w(0) <= NOT wire_Lshiftsmall_w_sel_w_range289w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range311w315w(0) <= NOT wire_Lshiftsmall_w_sel_w_range311w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range333w337w(0) <= NOT wire_Lshiftsmall_w_sel_w_range333w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range355w359w(0) <= NOT wire_Lshiftsmall_w_sel_w_range355w(0);
	loop15 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range268w280w281w282w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range268w280w281w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range268w276w277w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range289w301w302w303w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range289w301w302w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range289w297w298w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range311w323w324w325w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range311w323w324w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range311w319w320w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range333w345w346w347w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range333w345w346w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range333w341w342w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range355w367w368w369w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range355w367w368w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range355w363w364w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w283w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range268w280w281w282w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range268w272w273w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w304w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range289w301w302w303w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range289w293w294w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w326w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range311w323w324w325w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range311w315w316w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w348w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range333w345w346w347w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range333w337w338w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w370w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range355w367w368w369w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range355w359w360w(i);
	END GENERATE loop24;
	dir_w <= ( dir_pipe(0) & dir_w(3 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(191 DOWNTO 160);
	sbit_w <= ( sbit_piper1d & smux_w(127 DOWNTO 0) & data);
	sel_w <= ( distance(4 DOWNTO 0));
	smux_w <= ( wire_Lshiftsmall_w370w & wire_Lshiftsmall_w348w & wire_Lshiftsmall_w326w & wire_Lshiftsmall_w304w & wire_Lshiftsmall_w283w);
	wire_Lshiftsmall_w275w <= ( pad_w(0) & sbit_w(31 DOWNTO 1));
	wire_Lshiftsmall_w278w <= ( sbit_w(30 DOWNTO 0) & pad_w(0));
	wire_Lshiftsmall_w296w <= ( pad_w(1 DOWNTO 0) & sbit_w(63 DOWNTO 34));
	wire_Lshiftsmall_w299w <= ( sbit_w(61 DOWNTO 32) & pad_w(1 DOWNTO 0));
	wire_Lshiftsmall_w318w <= ( pad_w(3 DOWNTO 0) & sbit_w(95 DOWNTO 68));
	wire_Lshiftsmall_w321w <= ( sbit_w(91 DOWNTO 64) & pad_w(3 DOWNTO 0));
	wire_Lshiftsmall_w340w <= ( pad_w(7 DOWNTO 0) & sbit_w(127 DOWNTO 104));
	wire_Lshiftsmall_w343w <= ( sbit_w(119 DOWNTO 96) & pad_w(7 DOWNTO 0));
	wire_Lshiftsmall_w362w <= ( pad_w(15 DOWNTO 0) & sbit_w(159 DOWNTO 144));
	wire_Lshiftsmall_w365w <= ( sbit_w(143 DOWNTO 128) & pad_w(15 DOWNTO 0));
	wire_Lshiftsmall_w_dir_w_range265w(0) <= dir_w(0);
	wire_Lshiftsmall_w_dir_w_range287w(0) <= dir_w(1);
	wire_Lshiftsmall_w_dir_w_range308w(0) <= dir_w(2);
	wire_Lshiftsmall_w_dir_w_range330w(0) <= dir_w(3);
	wire_Lshiftsmall_w_dir_w_range352w(0) <= dir_w(4);
	wire_Lshiftsmall_w_sbit_w_range328w <= sbit_w(127 DOWNTO 96);
	wire_Lshiftsmall_w_sbit_w_range350w <= sbit_w(159 DOWNTO 128);
	wire_Lshiftsmall_w_sbit_w_range263w <= sbit_w(31 DOWNTO 0);
	wire_Lshiftsmall_w_sbit_w_range286w <= sbit_w(63 DOWNTO 32);
	wire_Lshiftsmall_w_sbit_w_range306w <= sbit_w(95 DOWNTO 64);
	wire_Lshiftsmall_w_sel_w_range268w(0) <= sel_w(0);
	wire_Lshiftsmall_w_sel_w_range289w(0) <= sel_w(1);
	wire_Lshiftsmall_w_sel_w_range311w(0) <= sel_w(2);
	wire_Lshiftsmall_w_sel_w_range333w(0) <= sel_w(3);
	wire_Lshiftsmall_w_sel_w_range355w(0) <= sel_w(4);
	wire_Lshiftsmall_w_smux_w_range371w <= smux_w(159 DOWNTO 128);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe(0) <= ( dir_w(4));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_Lshiftsmall_w_smux_w_range371w;
			END IF;
		END IF;
	END PROCESS;

 END RTL; --fplog_altbarrel_shift_itd


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" SHIFTDIR="LEFT" WIDTH=64 WIDTHDIST=6 data distance result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altbarrel_shift_qab IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (63 DOWNTO 0)
	 ); 
 END fplog_altbarrel_shift_qab;

 ARCHITECTURE RTL OF fplog_altbarrel_shift_qab IS

	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range382w394w395w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range382w390w391w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range403w415w416w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range403w411w412w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range425w437w438w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range425w433w434w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range447w459w460w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range447w455w456w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range469w481w482w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range469w477w478w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range491w503w504w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range491w499w500w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range382w386w387w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range403w407w408w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range425w429w430w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range447w451w452w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range469w473w474w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range491w495w496w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range382w394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range382w390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range403w415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range403w411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range425w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range425w433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range447w459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range447w455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range469w481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range469w477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range491w503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range491w499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range379w393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range401w414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range422w436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range444w458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range466w480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range488w502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range382w386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range403w407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range425w429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range447w451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range469w473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range491w495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range382w394w395w396w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range403w415w416w417w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range425w437w438w439w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range447w459w460w461w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range469w481w482w483w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range491w503w504w505w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w397w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w418w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w440w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w462w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w484w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w506w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (447 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (383 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w389w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w392w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w410w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w413w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w432w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w435w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w454w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w457w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w476w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w479w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w498w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w501w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range400w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range420w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range442w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range464w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range486w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range377w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	loop25 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range382w394w395w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range382w394w(0) AND wire_lzc_norm_L_w392w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range382w390w391w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range382w390w(0) AND wire_lzc_norm_L_w389w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range403w415w416w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range403w415w(0) AND wire_lzc_norm_L_w413w(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range403w411w412w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range403w411w(0) AND wire_lzc_norm_L_w410w(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range425w437w438w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range425w437w(0) AND wire_lzc_norm_L_w435w(i);
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range425w433w434w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range425w433w(0) AND wire_lzc_norm_L_w432w(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range447w459w460w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range447w459w(0) AND wire_lzc_norm_L_w457w(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range447w455w456w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range447w455w(0) AND wire_lzc_norm_L_w454w(i);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range469w481w482w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range469w481w(0) AND wire_lzc_norm_L_w479w(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range469w477w478w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range469w477w(0) AND wire_lzc_norm_L_w476w(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range491w503w504w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range491w503w(0) AND wire_lzc_norm_L_w501w(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range491w499w500w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range491w499w(0) AND wire_lzc_norm_L_w498w(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range382w386w387w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range382w386w(0) AND wire_lzc_norm_L_w_sbit_w_range377w(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range403w407w408w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range403w407w(0) AND wire_lzc_norm_L_w_sbit_w_range400w(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range425w429w430w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range425w429w(0) AND wire_lzc_norm_L_w_sbit_w_range420w(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range447w451w452w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range447w451w(0) AND wire_lzc_norm_L_w_sbit_w_range442w(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range469w473w474w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range469w473w(0) AND wire_lzc_norm_L_w_sbit_w_range464w(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range491w495w496w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range491w495w(0) AND wire_lzc_norm_L_w_sbit_w_range486w(i);
	END GENERATE loop42;
	wire_lzc_norm_L_w_lg_w_sel_w_range382w394w(0) <= wire_lzc_norm_L_w_sel_w_range382w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range379w393w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range382w390w(0) <= wire_lzc_norm_L_w_sel_w_range382w(0) AND wire_lzc_norm_L_w_dir_w_range379w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range403w415w(0) <= wire_lzc_norm_L_w_sel_w_range403w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range401w414w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range403w411w(0) <= wire_lzc_norm_L_w_sel_w_range403w(0) AND wire_lzc_norm_L_w_dir_w_range401w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range425w437w(0) <= wire_lzc_norm_L_w_sel_w_range425w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range422w436w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range425w433w(0) <= wire_lzc_norm_L_w_sel_w_range425w(0) AND wire_lzc_norm_L_w_dir_w_range422w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range447w459w(0) <= wire_lzc_norm_L_w_sel_w_range447w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range444w458w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range447w455w(0) <= wire_lzc_norm_L_w_sel_w_range447w(0) AND wire_lzc_norm_L_w_dir_w_range444w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range469w481w(0) <= wire_lzc_norm_L_w_sel_w_range469w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range466w480w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range469w477w(0) <= wire_lzc_norm_L_w_sel_w_range469w(0) AND wire_lzc_norm_L_w_dir_w_range466w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range491w503w(0) <= wire_lzc_norm_L_w_sel_w_range491w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range488w502w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range491w499w(0) <= wire_lzc_norm_L_w_sel_w_range491w(0) AND wire_lzc_norm_L_w_dir_w_range488w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range379w393w(0) <= NOT wire_lzc_norm_L_w_dir_w_range379w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range401w414w(0) <= NOT wire_lzc_norm_L_w_dir_w_range401w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range422w436w(0) <= NOT wire_lzc_norm_L_w_dir_w_range422w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range444w458w(0) <= NOT wire_lzc_norm_L_w_dir_w_range444w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range466w480w(0) <= NOT wire_lzc_norm_L_w_dir_w_range466w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range488w502w(0) <= NOT wire_lzc_norm_L_w_dir_w_range488w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range382w386w(0) <= NOT wire_lzc_norm_L_w_sel_w_range382w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range403w407w(0) <= NOT wire_lzc_norm_L_w_sel_w_range403w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range425w429w(0) <= NOT wire_lzc_norm_L_w_sel_w_range425w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range447w451w(0) <= NOT wire_lzc_norm_L_w_sel_w_range447w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range469w473w(0) <= NOT wire_lzc_norm_L_w_sel_w_range469w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range491w495w(0) <= NOT wire_lzc_norm_L_w_sel_w_range491w(0);
	loop43 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range382w394w395w396w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range382w394w395w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range382w390w391w(i);
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range403w415w416w417w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range403w415w416w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range403w411w412w(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range425w437w438w439w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range425w437w438w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range425w433w434w(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range447w459w460w461w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range447w459w460w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range447w455w456w(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range469w481w482w483w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range469w481w482w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range469w477w478w(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range491w503w504w505w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range491w503w504w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range491w499w500w(i);
	END GENERATE loop48;
	loop49 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w397w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range382w394w395w396w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range382w386w387w(i);
	END GENERATE loop49;
	loop50 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w418w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range403w415w416w417w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range403w407w408w(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w440w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range425w437w438w439w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range425w429w430w(i);
	END GENERATE loop51;
	loop52 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w462w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range447w459w460w461w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range447w451w452w(i);
	END GENERATE loop52;
	loop53 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w484w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range469w481w482w483w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range469w473w474w(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w506w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range491w503w504w505w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range491w495w496w(i);
	END GENERATE loop54;
	dir_w <= ( dir_w(5 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(447 DOWNTO 384);
	sbit_w <= ( smux_w(383 DOWNTO 0) & data);
	sel_w <= ( distance(5 DOWNTO 0));
	smux_w <= ( wire_lzc_norm_L_w506w & wire_lzc_norm_L_w484w & wire_lzc_norm_L_w462w & wire_lzc_norm_L_w440w & wire_lzc_norm_L_w418w & wire_lzc_norm_L_w397w);
	wire_lzc_norm_L_w389w <= ( pad_w(0) & sbit_w(63 DOWNTO 1));
	wire_lzc_norm_L_w392w <= ( sbit_w(62 DOWNTO 0) & pad_w(0));
	wire_lzc_norm_L_w410w <= ( pad_w(1 DOWNTO 0) & sbit_w(127 DOWNTO 66));
	wire_lzc_norm_L_w413w <= ( sbit_w(125 DOWNTO 64) & pad_w(1 DOWNTO 0));
	wire_lzc_norm_L_w432w <= ( pad_w(3 DOWNTO 0) & sbit_w(191 DOWNTO 132));
	wire_lzc_norm_L_w435w <= ( sbit_w(187 DOWNTO 128) & pad_w(3 DOWNTO 0));
	wire_lzc_norm_L_w454w <= ( pad_w(7 DOWNTO 0) & sbit_w(255 DOWNTO 200));
	wire_lzc_norm_L_w457w <= ( sbit_w(247 DOWNTO 192) & pad_w(7 DOWNTO 0));
	wire_lzc_norm_L_w476w <= ( pad_w(15 DOWNTO 0) & sbit_w(319 DOWNTO 272));
	wire_lzc_norm_L_w479w <= ( sbit_w(303 DOWNTO 256) & pad_w(15 DOWNTO 0));
	wire_lzc_norm_L_w498w <= ( pad_w(31 DOWNTO 0) & sbit_w(383 DOWNTO 352));
	wire_lzc_norm_L_w501w <= ( sbit_w(351 DOWNTO 320) & pad_w(31 DOWNTO 0));
	wire_lzc_norm_L_w_dir_w_range379w(0) <= dir_w(0);
	wire_lzc_norm_L_w_dir_w_range401w(0) <= dir_w(1);
	wire_lzc_norm_L_w_dir_w_range422w(0) <= dir_w(2);
	wire_lzc_norm_L_w_dir_w_range444w(0) <= dir_w(3);
	wire_lzc_norm_L_w_dir_w_range466w(0) <= dir_w(4);
	wire_lzc_norm_L_w_dir_w_range488w(0) <= dir_w(5);
	wire_lzc_norm_L_w_sbit_w_range400w <= sbit_w(127 DOWNTO 64);
	wire_lzc_norm_L_w_sbit_w_range420w <= sbit_w(191 DOWNTO 128);
	wire_lzc_norm_L_w_sbit_w_range442w <= sbit_w(255 DOWNTO 192);
	wire_lzc_norm_L_w_sbit_w_range464w <= sbit_w(319 DOWNTO 256);
	wire_lzc_norm_L_w_sbit_w_range486w <= sbit_w(383 DOWNTO 320);
	wire_lzc_norm_L_w_sbit_w_range377w <= sbit_w(63 DOWNTO 0);
	wire_lzc_norm_L_w_sel_w_range382w(0) <= sel_w(0);
	wire_lzc_norm_L_w_sel_w_range403w(0) <= sel_w(1);
	wire_lzc_norm_L_w_sel_w_range425w(0) <= sel_w(2);
	wire_lzc_norm_L_w_sel_w_range447w(0) <= sel_w(3);
	wire_lzc_norm_L_w_sel_w_range469w(0) <= sel_w(4);
	wire_lzc_norm_L_w_sel_w_range491w(0) <= sel_w(5);

 END RTL; --fplog_altbarrel_shift_qab


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" PIPELINE=1 SHIFTDIR="RIGHT" WIDTH=32 WIDTHDIST=5 aclr clk_en clock data distance result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END

--synthesis_resources = reg 33 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altbarrel_shift_51e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END fplog_altbarrel_shift_51e;

 ARCHITECTURE RTL OF fplog_altbarrel_shift_51e IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range518w530w531w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range518w526w527w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range539w551w552w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range539w547w548w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range561w573w574w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range561w569w570w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range583w595w596w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range583w591w592w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range605w617w618w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range605w613w614w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range518w522w523w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range539w543w544w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range561w565w566w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range583w587w588w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range605w609w610w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range518w530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range518w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range539w551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range539w547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range561w573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range561w569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range583w595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range583w591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range605w617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range605w613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_dir_w_range515w529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_dir_w_range537w550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_dir_w_range558w572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_dir_w_range580w594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_dir_w_range602w616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range518w522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range539w543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range561w565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range583w587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range605w609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range518w530w531w532w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range539w551w552w553w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range561w573w574w575w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range583w595w596w597w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range605w617w618w619w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w533w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w554w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w576w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w598w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w620w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (191 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (159 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w525w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w528w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w546w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w549w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w568w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w571w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w590w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w593w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w612w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w615w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_dir_w_range515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_dir_w_range537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_dir_w_range558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_dir_w_range580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_dir_w_range602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sbit_w_range578w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sbit_w_range600w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sbit_w_range513w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sbit_w_range536w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sbit_w_range556w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sel_w_range518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sel_w_range539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sel_w_range561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sel_w_range583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sel_w_range605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_smux_w_range621w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop55 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range518w530w531w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range518w530w(0) AND wire_Rshiftsmall_w528w(i);
	END GENERATE loop55;
	loop56 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range518w526w527w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range518w526w(0) AND wire_Rshiftsmall_w525w(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range539w551w552w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range539w551w(0) AND wire_Rshiftsmall_w549w(i);
	END GENERATE loop57;
	loop58 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range539w547w548w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range539w547w(0) AND wire_Rshiftsmall_w546w(i);
	END GENERATE loop58;
	loop59 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range561w573w574w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range561w573w(0) AND wire_Rshiftsmall_w571w(i);
	END GENERATE loop59;
	loop60 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range561w569w570w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range561w569w(0) AND wire_Rshiftsmall_w568w(i);
	END GENERATE loop60;
	loop61 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range583w595w596w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range583w595w(0) AND wire_Rshiftsmall_w593w(i);
	END GENERATE loop61;
	loop62 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range583w591w592w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range583w591w(0) AND wire_Rshiftsmall_w590w(i);
	END GENERATE loop62;
	loop63 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range605w617w618w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range605w617w(0) AND wire_Rshiftsmall_w615w(i);
	END GENERATE loop63;
	loop64 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range605w613w614w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range605w613w(0) AND wire_Rshiftsmall_w612w(i);
	END GENERATE loop64;
	loop65 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range518w522w523w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range518w522w(0) AND wire_Rshiftsmall_w_sbit_w_range513w(i);
	END GENERATE loop65;
	loop66 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range539w543w544w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range539w543w(0) AND wire_Rshiftsmall_w_sbit_w_range536w(i);
	END GENERATE loop66;
	loop67 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range561w565w566w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range561w565w(0) AND wire_Rshiftsmall_w_sbit_w_range556w(i);
	END GENERATE loop67;
	loop68 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range583w587w588w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range583w587w(0) AND wire_Rshiftsmall_w_sbit_w_range578w(i);
	END GENERATE loop68;
	loop69 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range605w609w610w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range605w609w(0) AND wire_Rshiftsmall_w_sbit_w_range600w(i);
	END GENERATE loop69;
	wire_Rshiftsmall_w_lg_w_sel_w_range518w530w(0) <= wire_Rshiftsmall_w_sel_w_range518w(0) AND wire_Rshiftsmall_w_lg_w_dir_w_range515w529w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range518w526w(0) <= wire_Rshiftsmall_w_sel_w_range518w(0) AND wire_Rshiftsmall_w_dir_w_range515w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range539w551w(0) <= wire_Rshiftsmall_w_sel_w_range539w(0) AND wire_Rshiftsmall_w_lg_w_dir_w_range537w550w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range539w547w(0) <= wire_Rshiftsmall_w_sel_w_range539w(0) AND wire_Rshiftsmall_w_dir_w_range537w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range561w573w(0) <= wire_Rshiftsmall_w_sel_w_range561w(0) AND wire_Rshiftsmall_w_lg_w_dir_w_range558w572w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range561w569w(0) <= wire_Rshiftsmall_w_sel_w_range561w(0) AND wire_Rshiftsmall_w_dir_w_range558w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range583w595w(0) <= wire_Rshiftsmall_w_sel_w_range583w(0) AND wire_Rshiftsmall_w_lg_w_dir_w_range580w594w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range583w591w(0) <= wire_Rshiftsmall_w_sel_w_range583w(0) AND wire_Rshiftsmall_w_dir_w_range580w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range605w617w(0) <= wire_Rshiftsmall_w_sel_w_range605w(0) AND wire_Rshiftsmall_w_lg_w_dir_w_range602w616w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range605w613w(0) <= wire_Rshiftsmall_w_sel_w_range605w(0) AND wire_Rshiftsmall_w_dir_w_range602w(0);
	wire_Rshiftsmall_w_lg_w_dir_w_range515w529w(0) <= NOT wire_Rshiftsmall_w_dir_w_range515w(0);
	wire_Rshiftsmall_w_lg_w_dir_w_range537w550w(0) <= NOT wire_Rshiftsmall_w_dir_w_range537w(0);
	wire_Rshiftsmall_w_lg_w_dir_w_range558w572w(0) <= NOT wire_Rshiftsmall_w_dir_w_range558w(0);
	wire_Rshiftsmall_w_lg_w_dir_w_range580w594w(0) <= NOT wire_Rshiftsmall_w_dir_w_range580w(0);
	wire_Rshiftsmall_w_lg_w_dir_w_range602w616w(0) <= NOT wire_Rshiftsmall_w_dir_w_range602w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range518w522w(0) <= NOT wire_Rshiftsmall_w_sel_w_range518w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range539w543w(0) <= NOT wire_Rshiftsmall_w_sel_w_range539w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range561w565w(0) <= NOT wire_Rshiftsmall_w_sel_w_range561w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range583w587w(0) <= NOT wire_Rshiftsmall_w_sel_w_range583w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range605w609w(0) <= NOT wire_Rshiftsmall_w_sel_w_range605w(0);
	loop70 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range518w530w531w532w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range518w530w531w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range518w526w527w(i);
	END GENERATE loop70;
	loop71 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range539w551w552w553w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range539w551w552w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range539w547w548w(i);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range561w573w574w575w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range561w573w574w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range561w569w570w(i);
	END GENERATE loop72;
	loop73 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range583w595w596w597w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range583w595w596w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range583w591w592w(i);
	END GENERATE loop73;
	loop74 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range605w617w618w619w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range605w617w618w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range605w613w614w(i);
	END GENERATE loop74;
	loop75 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w533w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range518w530w531w532w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range518w522w523w(i);
	END GENERATE loop75;
	loop76 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w554w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range539w551w552w553w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range539w543w544w(i);
	END GENERATE loop76;
	loop77 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w576w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range561w573w574w575w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range561w565w566w(i);
	END GENERATE loop77;
	loop78 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w598w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range583w595w596w597w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range583w587w588w(i);
	END GENERATE loop78;
	loop79 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w620w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range605w617w618w619w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range605w609w610w(i);
	END GENERATE loop79;
	dir_w <= ( dir_pipe(0) & dir_w(3 DOWNTO 0) & direction_w);
	direction_w <= '1';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(191 DOWNTO 160);
	sbit_w <= ( sbit_piper1d & smux_w(127 DOWNTO 0) & data);
	sel_w <= ( distance(4 DOWNTO 0));
	smux_w <= ( wire_Rshiftsmall_w620w & wire_Rshiftsmall_w598w & wire_Rshiftsmall_w576w & wire_Rshiftsmall_w554w & wire_Rshiftsmall_w533w);
	wire_Rshiftsmall_w525w <= ( pad_w(0) & sbit_w(31 DOWNTO 1));
	wire_Rshiftsmall_w528w <= ( sbit_w(30 DOWNTO 0) & pad_w(0));
	wire_Rshiftsmall_w546w <= ( pad_w(1 DOWNTO 0) & sbit_w(63 DOWNTO 34));
	wire_Rshiftsmall_w549w <= ( sbit_w(61 DOWNTO 32) & pad_w(1 DOWNTO 0));
	wire_Rshiftsmall_w568w <= ( pad_w(3 DOWNTO 0) & sbit_w(95 DOWNTO 68));
	wire_Rshiftsmall_w571w <= ( sbit_w(91 DOWNTO 64) & pad_w(3 DOWNTO 0));
	wire_Rshiftsmall_w590w <= ( pad_w(7 DOWNTO 0) & sbit_w(127 DOWNTO 104));
	wire_Rshiftsmall_w593w <= ( sbit_w(119 DOWNTO 96) & pad_w(7 DOWNTO 0));
	wire_Rshiftsmall_w612w <= ( pad_w(15 DOWNTO 0) & sbit_w(159 DOWNTO 144));
	wire_Rshiftsmall_w615w <= ( sbit_w(143 DOWNTO 128) & pad_w(15 DOWNTO 0));
	wire_Rshiftsmall_w_dir_w_range515w(0) <= dir_w(0);
	wire_Rshiftsmall_w_dir_w_range537w(0) <= dir_w(1);
	wire_Rshiftsmall_w_dir_w_range558w(0) <= dir_w(2);
	wire_Rshiftsmall_w_dir_w_range580w(0) <= dir_w(3);
	wire_Rshiftsmall_w_dir_w_range602w(0) <= dir_w(4);
	wire_Rshiftsmall_w_sbit_w_range578w <= sbit_w(127 DOWNTO 96);
	wire_Rshiftsmall_w_sbit_w_range600w <= sbit_w(159 DOWNTO 128);
	wire_Rshiftsmall_w_sbit_w_range513w <= sbit_w(31 DOWNTO 0);
	wire_Rshiftsmall_w_sbit_w_range536w <= sbit_w(63 DOWNTO 32);
	wire_Rshiftsmall_w_sbit_w_range556w <= sbit_w(95 DOWNTO 64);
	wire_Rshiftsmall_w_sel_w_range518w(0) <= sel_w(0);
	wire_Rshiftsmall_w_sel_w_range539w(0) <= sel_w(1);
	wire_Rshiftsmall_w_sel_w_range561w(0) <= sel_w(2);
	wire_Rshiftsmall_w_sel_w_range583w(0) <= sel_w(3);
	wire_Rshiftsmall_w_sel_w_range605w(0) <= sel_w(4);
	wire_Rshiftsmall_w_smux_w_range621w <= smux_w(159 DOWNTO 128);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe(0) <= ( dir_w(4));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_Rshiftsmall_w_smux_w_range621w;
			END IF;
		END IF;
	END PROCESS;

 END RTL; --fplog_altbarrel_shift_51e


--altfp_log_and_or CBX_AUTO_BLACKBOX="ALL" LUT_INPUT_COUNT=6 OPERATION="AND" PIPELINE=3 WIDTH=8 aclr clken clock data result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

--synthesis_resources = reg 4 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_and_or_h9b IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC
	 ); 
 END fplog_altfp_log_and_or_h9b;

 ARCHITECTURE RTL OF fplog_altfp_log_and_or_h9b IS

	 SIGNAL	 connection_dffe0	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range628w632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range631w635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range634w638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range637w641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range640w644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range646w649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r2_w_range655w659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  connection_r0_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  connection_r1_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  connection_r2_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  operation_r1_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  operation_r2_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r1_w_range657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r2_w_range655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_exp_nan_w_lg_w_operation_r1_w_range628w632w(0) <= wire_exp_nan_w_operation_r1_w_range628w(0) AND wire_exp_nan_w_connection_r0_w_range630w(0);
	wire_exp_nan_w_lg_w_operation_r1_w_range631w635w(0) <= wire_exp_nan_w_operation_r1_w_range631w(0) AND wire_exp_nan_w_connection_r0_w_range633w(0);
	wire_exp_nan_w_lg_w_operation_r1_w_range634w638w(0) <= wire_exp_nan_w_operation_r1_w_range634w(0) AND wire_exp_nan_w_connection_r0_w_range636w(0);
	wire_exp_nan_w_lg_w_operation_r1_w_range637w641w(0) <= wire_exp_nan_w_operation_r1_w_range637w(0) AND wire_exp_nan_w_connection_r0_w_range639w(0);
	wire_exp_nan_w_lg_w_operation_r1_w_range640w644w(0) <= wire_exp_nan_w_operation_r1_w_range640w(0) AND wire_exp_nan_w_connection_r0_w_range642w(0);
	wire_exp_nan_w_lg_w_operation_r1_w_range646w649w(0) <= wire_exp_nan_w_operation_r1_w_range646w(0) AND wire_exp_nan_w_connection_r0_w_range647w(0);
	wire_exp_nan_w_lg_w_operation_r2_w_range655w659w(0) <= wire_exp_nan_w_operation_r2_w_range655w(0) AND wire_exp_nan_w_connection_r1_w_range657w(0);
	connection_r0_w <= data;
	connection_r1_w <= connection_dffe0;
	connection_r2_w <= connection_dffe1;
	operation_r1_w <= ( wire_exp_nan_w_lg_w_operation_r1_w_range646w649w & connection_r0_w(6) & wire_exp_nan_w_lg_w_operation_r1_w_range640w644w & wire_exp_nan_w_lg_w_operation_r1_w_range637w641w & wire_exp_nan_w_lg_w_operation_r1_w_range634w638w & wire_exp_nan_w_lg_w_operation_r1_w_range631w635w & wire_exp_nan_w_lg_w_operation_r1_w_range628w632w & connection_r0_w(0));
	operation_r2_w <= ( wire_exp_nan_w_lg_w_operation_r2_w_range655w659w & connection_r1_w(0));
	result <= connection_dffe2;
	wire_exp_nan_w_connection_r0_w_range630w(0) <= connection_r0_w(1);
	wire_exp_nan_w_connection_r0_w_range633w(0) <= connection_r0_w(2);
	wire_exp_nan_w_connection_r0_w_range636w(0) <= connection_r0_w(3);
	wire_exp_nan_w_connection_r0_w_range639w(0) <= connection_r0_w(4);
	wire_exp_nan_w_connection_r0_w_range642w(0) <= connection_r0_w(5);
	wire_exp_nan_w_connection_r0_w_range647w(0) <= connection_r0_w(7);
	wire_exp_nan_w_connection_r1_w_range657w(0) <= connection_r1_w(1);
	wire_exp_nan_w_operation_r1_w_range628w(0) <= operation_r1_w(0);
	wire_exp_nan_w_operation_r1_w_range631w(0) <= operation_r1_w(1);
	wire_exp_nan_w_operation_r1_w_range634w(0) <= operation_r1_w(2);
	wire_exp_nan_w_operation_r1_w_range637w(0) <= operation_r1_w(3);
	wire_exp_nan_w_operation_r1_w_range640w(0) <= operation_r1_w(4);
	wire_exp_nan_w_operation_r1_w_range646w(0) <= operation_r1_w(6);
	wire_exp_nan_w_operation_r2_w_range655w(0) <= operation_r2_w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe0 <= ( operation_r1_w(7) & operation_r1_w(5));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe1(0) <= ( operation_r2_w(1));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe2 <= connection_r2_w(0);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --fplog_altfp_log_and_or_h9b


--altfp_log_and_or CBX_AUTO_BLACKBOX="ALL" LUT_INPUT_COUNT=6 OPERATION="OR" PIPELINE=3 WIDTH=8 aclr clken clock data result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

--synthesis_resources = reg 4 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_and_or_v6b IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC
	 ); 
 END fplog_altfp_log_and_or_v6b;

 ARCHITECTURE RTL OF fplog_altfp_log_and_or_v6b IS

	 SIGNAL	 connection_dffe0	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range664w668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range667w671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range670w674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range673w677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range676w680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range682w685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r2_w_range691w695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  connection_r0_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  connection_r1_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  connection_r2_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  operation_r1_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  operation_r2_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r1_w_range693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r2_w_range691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_exp_zero_w_lg_w_operation_r1_w_range664w668w(0) <= wire_exp_zero_w_operation_r1_w_range664w(0) OR wire_exp_zero_w_connection_r0_w_range666w(0);
	wire_exp_zero_w_lg_w_operation_r1_w_range667w671w(0) <= wire_exp_zero_w_operation_r1_w_range667w(0) OR wire_exp_zero_w_connection_r0_w_range669w(0);
	wire_exp_zero_w_lg_w_operation_r1_w_range670w674w(0) <= wire_exp_zero_w_operation_r1_w_range670w(0) OR wire_exp_zero_w_connection_r0_w_range672w(0);
	wire_exp_zero_w_lg_w_operation_r1_w_range673w677w(0) <= wire_exp_zero_w_operation_r1_w_range673w(0) OR wire_exp_zero_w_connection_r0_w_range675w(0);
	wire_exp_zero_w_lg_w_operation_r1_w_range676w680w(0) <= wire_exp_zero_w_operation_r1_w_range676w(0) OR wire_exp_zero_w_connection_r0_w_range678w(0);
	wire_exp_zero_w_lg_w_operation_r1_w_range682w685w(0) <= wire_exp_zero_w_operation_r1_w_range682w(0) OR wire_exp_zero_w_connection_r0_w_range683w(0);
	wire_exp_zero_w_lg_w_operation_r2_w_range691w695w(0) <= wire_exp_zero_w_operation_r2_w_range691w(0) OR wire_exp_zero_w_connection_r1_w_range693w(0);
	connection_r0_w <= data;
	connection_r1_w <= connection_dffe0;
	connection_r2_w <= connection_dffe1;
	operation_r1_w <= ( wire_exp_zero_w_lg_w_operation_r1_w_range682w685w & connection_r0_w(6) & wire_exp_zero_w_lg_w_operation_r1_w_range676w680w & wire_exp_zero_w_lg_w_operation_r1_w_range673w677w & wire_exp_zero_w_lg_w_operation_r1_w_range670w674w & wire_exp_zero_w_lg_w_operation_r1_w_range667w671w & wire_exp_zero_w_lg_w_operation_r1_w_range664w668w & connection_r0_w(0));
	operation_r2_w <= ( wire_exp_zero_w_lg_w_operation_r2_w_range691w695w & connection_r1_w(0));
	result <= connection_dffe2;
	wire_exp_zero_w_connection_r0_w_range666w(0) <= connection_r0_w(1);
	wire_exp_zero_w_connection_r0_w_range669w(0) <= connection_r0_w(2);
	wire_exp_zero_w_connection_r0_w_range672w(0) <= connection_r0_w(3);
	wire_exp_zero_w_connection_r0_w_range675w(0) <= connection_r0_w(4);
	wire_exp_zero_w_connection_r0_w_range678w(0) <= connection_r0_w(5);
	wire_exp_zero_w_connection_r0_w_range683w(0) <= connection_r0_w(7);
	wire_exp_zero_w_connection_r1_w_range693w(0) <= connection_r1_w(1);
	wire_exp_zero_w_operation_r1_w_range664w(0) <= operation_r1_w(0);
	wire_exp_zero_w_operation_r1_w_range667w(0) <= operation_r1_w(1);
	wire_exp_zero_w_operation_r1_w_range670w(0) <= operation_r1_w(2);
	wire_exp_zero_w_operation_r1_w_range673w(0) <= operation_r1_w(3);
	wire_exp_zero_w_operation_r1_w_range676w(0) <= operation_r1_w(4);
	wire_exp_zero_w_operation_r1_w_range682w(0) <= operation_r1_w(6);
	wire_exp_zero_w_operation_r2_w_range691w(0) <= operation_r2_w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe0 <= ( operation_r1_w(7) & operation_r1_w(5));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe1(0) <= ( operation_r2_w(1));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe2 <= connection_r2_w(0);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --fplog_altfp_log_and_or_v6b


--altfp_log_and_or CBX_AUTO_BLACKBOX="ALL" LUT_INPUT_COUNT=6 OPERATION="OR" PIPELINE=3 WIDTH=23 aclr clken clock data result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

--synthesis_resources = reg 6 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_and_or_c8b IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (22 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC
	 ); 
 END fplog_altfp_log_and_or_c8b;

 ARCHITECTURE RTL OF fplog_altfp_log_and_or_c8b IS

	 SIGNAL	 connection_dffe0	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range700w704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range729w733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range735w738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range737w741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range740w744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range743w747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range746w750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range752w755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range754w758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range703w707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range757w761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range760w764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range706w710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range709w713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range712w716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range718w721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range720w724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range723w727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range726w730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r2_w_range772w776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r2_w_range775w779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r2_w_range778w782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  connection_r0_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  connection_r1_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  connection_r2_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  operation_r1_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  operation_r2_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r1_w_range774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r1_w_range777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r1_w_range780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r2_w_range772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r2_w_range775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r2_w_range778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_man_inf_w_lg_w_operation_r1_w_range700w704w(0) <= wire_man_inf_w_operation_r1_w_range700w(0) OR wire_man_inf_w_connection_r0_w_range702w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range729w733w(0) <= wire_man_inf_w_operation_r1_w_range729w(0) OR wire_man_inf_w_connection_r0_w_range731w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range735w738w(0) <= wire_man_inf_w_operation_r1_w_range735w(0) OR wire_man_inf_w_connection_r0_w_range736w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range737w741w(0) <= wire_man_inf_w_operation_r1_w_range737w(0) OR wire_man_inf_w_connection_r0_w_range739w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range740w744w(0) <= wire_man_inf_w_operation_r1_w_range740w(0) OR wire_man_inf_w_connection_r0_w_range742w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range743w747w(0) <= wire_man_inf_w_operation_r1_w_range743w(0) OR wire_man_inf_w_connection_r0_w_range745w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range746w750w(0) <= wire_man_inf_w_operation_r1_w_range746w(0) OR wire_man_inf_w_connection_r0_w_range748w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range752w755w(0) <= wire_man_inf_w_operation_r1_w_range752w(0) OR wire_man_inf_w_connection_r0_w_range753w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range754w758w(0) <= wire_man_inf_w_operation_r1_w_range754w(0) OR wire_man_inf_w_connection_r0_w_range756w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range703w707w(0) <= wire_man_inf_w_operation_r1_w_range703w(0) OR wire_man_inf_w_connection_r0_w_range705w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range757w761w(0) <= wire_man_inf_w_operation_r1_w_range757w(0) OR wire_man_inf_w_connection_r0_w_range759w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range760w764w(0) <= wire_man_inf_w_operation_r1_w_range760w(0) OR wire_man_inf_w_connection_r0_w_range762w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range706w710w(0) <= wire_man_inf_w_operation_r1_w_range706w(0) OR wire_man_inf_w_connection_r0_w_range708w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range709w713w(0) <= wire_man_inf_w_operation_r1_w_range709w(0) OR wire_man_inf_w_connection_r0_w_range711w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range712w716w(0) <= wire_man_inf_w_operation_r1_w_range712w(0) OR wire_man_inf_w_connection_r0_w_range714w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range718w721w(0) <= wire_man_inf_w_operation_r1_w_range718w(0) OR wire_man_inf_w_connection_r0_w_range719w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range720w724w(0) <= wire_man_inf_w_operation_r1_w_range720w(0) OR wire_man_inf_w_connection_r0_w_range722w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range723w727w(0) <= wire_man_inf_w_operation_r1_w_range723w(0) OR wire_man_inf_w_connection_r0_w_range725w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range726w730w(0) <= wire_man_inf_w_operation_r1_w_range726w(0) OR wire_man_inf_w_connection_r0_w_range728w(0);
	wire_man_inf_w_lg_w_operation_r2_w_range772w776w(0) <= wire_man_inf_w_operation_r2_w_range772w(0) OR wire_man_inf_w_connection_r1_w_range774w(0);
	wire_man_inf_w_lg_w_operation_r2_w_range775w779w(0) <= wire_man_inf_w_operation_r2_w_range775w(0) OR wire_man_inf_w_connection_r1_w_range777w(0);
	wire_man_inf_w_lg_w_operation_r2_w_range778w782w(0) <= wire_man_inf_w_operation_r2_w_range778w(0) OR wire_man_inf_w_connection_r1_w_range780w(0);
	connection_r0_w <= data;
	connection_r1_w <= connection_dffe0;
	connection_r2_w <= connection_dffe1;
	operation_r1_w <= ( wire_man_inf_w_lg_w_operation_r1_w_range760w764w & wire_man_inf_w_lg_w_operation_r1_w_range757w761w & wire_man_inf_w_lg_w_operation_r1_w_range754w758w & wire_man_inf_w_lg_w_operation_r1_w_range752w755w & connection_r0_w(18) & wire_man_inf_w_lg_w_operation_r1_w_range746w750w & wire_man_inf_w_lg_w_operation_r1_w_range743w747w & wire_man_inf_w_lg_w_operation_r1_w_range740w744w & wire_man_inf_w_lg_w_operation_r1_w_range737w741w & wire_man_inf_w_lg_w_operation_r1_w_range735w738w & connection_r0_w(12) & wire_man_inf_w_lg_w_operation_r1_w_range729w733w & wire_man_inf_w_lg_w_operation_r1_w_range726w730w & wire_man_inf_w_lg_w_operation_r1_w_range723w727w & wire_man_inf_w_lg_w_operation_r1_w_range720w724w & wire_man_inf_w_lg_w_operation_r1_w_range718w721w & connection_r0_w(6) & wire_man_inf_w_lg_w_operation_r1_w_range712w716w & wire_man_inf_w_lg_w_operation_r1_w_range709w713w & wire_man_inf_w_lg_w_operation_r1_w_range706w710w & wire_man_inf_w_lg_w_operation_r1_w_range703w707w & wire_man_inf_w_lg_w_operation_r1_w_range700w704w & connection_r0_w(0));
	operation_r2_w <= ( wire_man_inf_w_lg_w_operation_r2_w_range778w782w & wire_man_inf_w_lg_w_operation_r2_w_range775w779w & wire_man_inf_w_lg_w_operation_r2_w_range772w776w & connection_r1_w(0));
	result <= connection_dffe2;
	wire_man_inf_w_connection_r0_w_range728w(0) <= connection_r0_w(10);
	wire_man_inf_w_connection_r0_w_range731w(0) <= connection_r0_w(11);
	wire_man_inf_w_connection_r0_w_range736w(0) <= connection_r0_w(13);
	wire_man_inf_w_connection_r0_w_range739w(0) <= connection_r0_w(14);
	wire_man_inf_w_connection_r0_w_range742w(0) <= connection_r0_w(15);
	wire_man_inf_w_connection_r0_w_range745w(0) <= connection_r0_w(16);
	wire_man_inf_w_connection_r0_w_range748w(0) <= connection_r0_w(17);
	wire_man_inf_w_connection_r0_w_range753w(0) <= connection_r0_w(19);
	wire_man_inf_w_connection_r0_w_range702w(0) <= connection_r0_w(1);
	wire_man_inf_w_connection_r0_w_range756w(0) <= connection_r0_w(20);
	wire_man_inf_w_connection_r0_w_range759w(0) <= connection_r0_w(21);
	wire_man_inf_w_connection_r0_w_range762w(0) <= connection_r0_w(22);
	wire_man_inf_w_connection_r0_w_range705w(0) <= connection_r0_w(2);
	wire_man_inf_w_connection_r0_w_range708w(0) <= connection_r0_w(3);
	wire_man_inf_w_connection_r0_w_range711w(0) <= connection_r0_w(4);
	wire_man_inf_w_connection_r0_w_range714w(0) <= connection_r0_w(5);
	wire_man_inf_w_connection_r0_w_range719w(0) <= connection_r0_w(7);
	wire_man_inf_w_connection_r0_w_range722w(0) <= connection_r0_w(8);
	wire_man_inf_w_connection_r0_w_range725w(0) <= connection_r0_w(9);
	wire_man_inf_w_connection_r1_w_range774w(0) <= connection_r1_w(1);
	wire_man_inf_w_connection_r1_w_range777w(0) <= connection_r1_w(2);
	wire_man_inf_w_connection_r1_w_range780w(0) <= connection_r1_w(3);
	wire_man_inf_w_operation_r1_w_range700w(0) <= operation_r1_w(0);
	wire_man_inf_w_operation_r1_w_range729w(0) <= operation_r1_w(10);
	wire_man_inf_w_operation_r1_w_range735w(0) <= operation_r1_w(12);
	wire_man_inf_w_operation_r1_w_range737w(0) <= operation_r1_w(13);
	wire_man_inf_w_operation_r1_w_range740w(0) <= operation_r1_w(14);
	wire_man_inf_w_operation_r1_w_range743w(0) <= operation_r1_w(15);
	wire_man_inf_w_operation_r1_w_range746w(0) <= operation_r1_w(16);
	wire_man_inf_w_operation_r1_w_range752w(0) <= operation_r1_w(18);
	wire_man_inf_w_operation_r1_w_range754w(0) <= operation_r1_w(19);
	wire_man_inf_w_operation_r1_w_range703w(0) <= operation_r1_w(1);
	wire_man_inf_w_operation_r1_w_range757w(0) <= operation_r1_w(20);
	wire_man_inf_w_operation_r1_w_range760w(0) <= operation_r1_w(21);
	wire_man_inf_w_operation_r1_w_range706w(0) <= operation_r1_w(2);
	wire_man_inf_w_operation_r1_w_range709w(0) <= operation_r1_w(3);
	wire_man_inf_w_operation_r1_w_range712w(0) <= operation_r1_w(4);
	wire_man_inf_w_operation_r1_w_range718w(0) <= operation_r1_w(6);
	wire_man_inf_w_operation_r1_w_range720w(0) <= operation_r1_w(7);
	wire_man_inf_w_operation_r1_w_range723w(0) <= operation_r1_w(8);
	wire_man_inf_w_operation_r1_w_range726w(0) <= operation_r1_w(9);
	wire_man_inf_w_operation_r2_w_range772w(0) <= operation_r2_w(0);
	wire_man_inf_w_operation_r2_w_range775w(0) <= operation_r2_w(1);
	wire_man_inf_w_operation_r2_w_range778w(0) <= operation_r2_w(2);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe0 <= ( operation_r1_w(22) & operation_r1_w(17) & operation_r1_w(11) & operation_r1_w(5));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe1(0) <= ( operation_r2_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe2 <= connection_r2_w(0);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --fplog_altfp_log_and_or_c8b


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="ADD" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=39 aclr clken clock dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_s0e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (38 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (38 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (38 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_s0e;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_s0e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout793w794w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout792w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout793w794w795w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout793w794w795w & wire_csa_lower_result);
	loop80 : FOR i IN 0 TO 18 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout793w794w(i) <= wire_csa_lower_w_lg_cout793w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop80;
	loop81 : FOR i IN 0 TO 18 GENERATE 
		wire_csa_lower_w_lg_cout792w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop81;
	wire_csa_lower_w_lg_cout793w(0) <= NOT wire_csa_lower_cout;
	loop82 : FOR i IN 0 TO 18 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout793w794w795w(i) <= wire_csa_lower_w_lg_w_lg_cout793w794w(i) OR wire_csa_lower_w_lg_cout792w(i);
	END GENERATE loop82;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 20
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(19 DOWNTO 0),
		datab => datab(19 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 19
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(38 DOWNTO 20),
		datab => datab(38 DOWNTO 20),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 19
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(38 DOWNTO 20),
		datab => datab(38 DOWNTO 20),
		result => wire_csa_upper1_result
	  );

 END RTL; --fplog_altfp_log_csa_s0e


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="ADD" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=31 aclr clken clock dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_k0e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (30 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (30 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (30 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_k0e;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_k0e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout804w805w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout803w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout804w805w806w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout804w805w806w & wire_csa_lower_result);
	loop83 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout804w805w(i) <= wire_csa_lower_w_lg_cout804w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop83;
	loop84 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_cout803w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop84;
	wire_csa_lower_w_lg_cout804w(0) <= NOT wire_csa_lower_cout;
	loop85 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout804w805w806w(i) <= wire_csa_lower_w_lg_w_lg_cout804w805w(i) OR wire_csa_lower_w_lg_cout803w(i);
	END GENERATE loop85;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 16
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(15 DOWNTO 0),
		datab => datab(15 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(30 DOWNTO 16),
		datab => datab(30 DOWNTO 16),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(30 DOWNTO 16),
		datab => datab(30 DOWNTO 16),
		result => wire_csa_upper1_result
	  );

 END RTL; --fplog_altfp_log_csa_k0e


--altfp_log_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=8 dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_0nc IS 
	 PORT 
	 ( 
		 dataa	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_0nc;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_0nc IS

	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub1_result;
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		dataa => dataa,
		datab => datab,
		result => wire_add_sub1_result
	  );

 END RTL; --fplog_altfp_log_csa_0nc


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=12 dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_d4b IS 
	 PORT 
	 ( 
		 dataa	:	IN  STD_LOGIC_VECTOR (11 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (11 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (11 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_d4b;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_d4b IS

	 SIGNAL  wire_add_sub2_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub2_result;
	add_sub2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		dataa => dataa,
		datab => datab,
		result => wire_add_sub2_result
	  );

 END RTL; --fplog_altfp_log_csa_d4b


--altfp_log_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=6 dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_umc IS 
	 PORT 
	 ( 
		 dataa	:	IN  STD_LOGIC_VECTOR (5 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (5 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_umc;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_umc IS

	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub3_result;
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		dataa => dataa,
		datab => datab,
		result => wire_add_sub3_result
	  );

 END RTL; --fplog_altfp_log_csa_umc


--altfp_log_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=26 aclr clken clock dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_nlf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (25 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_nlf;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_nlf IS

	 SIGNAL  wire_add_sub4_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub4_result;
	add_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 26
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => wire_add_sub4_result
	  );

 END RTL; --fplog_altfp_log_csa_nlf


--altfp_log_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_PIPELINE=2 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=8 aclr clken clock dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_8kf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_8kf;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_8kf IS

	 SIGNAL  wire_add_sub5_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub5_result;
	add_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => wire_add_sub5_result
	  );

 END RTL; --fplog_altfp_log_csa_8kf


--altfp_log_rr_block CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" WIDTH_ALMOSTLOG=39 WIDTH_Y0=25 WIDTH_Z=26 a0_in aclr almostlog clk_en clock y0_in z
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="ADD" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=29 aclr clken clock dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_r0e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (28 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (28 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (28 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_r0e;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_r0e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout1193w1194w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1192w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout1193w1194w1195w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout1193w1194w1195w & wire_csa_lower_result);
	loop86 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout1193w1194w(i) <= wire_csa_lower_w_lg_cout1193w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop86;
	loop87 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_cout1192w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop87;
	wire_csa_lower_w_lg_cout1193w(0) <= NOT wire_csa_lower_cout;
	loop88 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout1193w1194w1195w(i) <= wire_csa_lower_w_lg_w_lg_cout1193w1194w(i) OR wire_csa_lower_w_lg_cout1192w(i);
	END GENERATE loop88;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(14 DOWNTO 0),
		datab => datab(14 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(28 DOWNTO 15),
		datab => datab(28 DOWNTO 15),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(28 DOWNTO 15),
		datab => datab(28 DOWNTO 15),
		result => wire_csa_upper1_result
	  );

 END RTL; --fplog_altfp_log_csa_r0e


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="ADD" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=26 aclr clken clock dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_o0e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (25 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_o0e;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_o0e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout1204w1205w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1203w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout1204w1205w1206w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout1204w1205w1206w & wire_csa_lower_result);
	loop89 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout1204w1205w(i) <= wire_csa_lower_w_lg_cout1204w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop89;
	loop90 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_cout1203w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop90;
	wire_csa_lower_w_lg_cout1204w(0) <= NOT wire_csa_lower_cout;
	loop91 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout1204w1205w1206w(i) <= wire_csa_lower_w_lg_w_lg_cout1204w1205w(i) OR wire_csa_lower_w_lg_cout1203w(i);
	END GENERATE loop91;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(12 DOWNTO 0),
		datab => datab(12 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(25 DOWNTO 13),
		datab => datab(25 DOWNTO 13),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(25 DOWNTO 13),
		datab => datab(25 DOWNTO 13),
		result => wire_csa_upper1_result
	  );

 END RTL; --fplog_altfp_log_csa_o0e


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=31 aclr clken clock dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_l1e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (30 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (30 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (30 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_l1e;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_l1e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout1215w1216w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1214w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout1215w1216w1217w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout1215w1216w1217w & wire_csa_lower_result);
	loop92 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout1215w1216w(i) <= wire_csa_lower_w_lg_cout1215w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop92;
	loop93 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_cout1214w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop93;
	wire_csa_lower_w_lg_cout1215w(0) <= NOT wire_csa_lower_cout;
	loop94 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout1215w1216w1217w(i) <= wire_csa_lower_w_lg_w_lg_cout1215w1216w(i) OR wire_csa_lower_w_lg_cout1214w(i);
	END GENERATE loop94;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 16
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(15 DOWNTO 0),
		datab => datab(15 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(30 DOWNTO 16),
		datab => datab(30 DOWNTO 16),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(30 DOWNTO 16),
		datab => datab(30 DOWNTO 16),
		result => wire_csa_upper1_result
	  );

 END RTL; --fplog_altfp_log_csa_l1e


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=29 aclr clken clock dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_s1e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (28 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (28 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (28 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_s1e;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_s1e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout1226w1227w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1225w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout1226w1227w1228w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout1226w1227w1228w & wire_csa_lower_result);
	loop95 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout1226w1227w(i) <= wire_csa_lower_w_lg_cout1226w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop95;
	loop96 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_cout1225w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop96;
	wire_csa_lower_w_lg_cout1226w(0) <= NOT wire_csa_lower_cout;
	loop97 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout1226w1227w1228w(i) <= wire_csa_lower_w_lg_w_lg_cout1226w1227w(i) OR wire_csa_lower_w_lg_cout1225w(i);
	END GENERATE loop97;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(14 DOWNTO 0),
		datab => datab(14 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(28 DOWNTO 15),
		datab => datab(28 DOWNTO 15),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(28 DOWNTO 15),
		datab => datab(28 DOWNTO 15),
		result => wire_csa_upper1_result
	  );

 END RTL; --fplog_altfp_log_csa_s1e


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=26 aclr clken clock dataa datab result
--VERSION_BEGIN 16.1 cbx_altbarrel_shift 2016:10:24:15:04:16:SJ cbx_altfp_log 2016:10:24:15:04:16:SJ cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_altsquare 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_mult 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_padd 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_csa_p1e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (25 DOWNTO 0)
	 ); 
 END fplog_altfp_log_csa_p1e;

 ARCHITECTURE RTL OF fplog_altfp_log_csa_p1e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout1237w1238w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1236w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout1237w1238w1239w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout1237w1238w1239w & wire_csa_lower_result);
	loop98 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout1237w1238w(i) <= wire_csa_lower_w_lg_cout1237w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop98;
	loop99 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_cout1236w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop99;
	wire_csa_lower_w_lg_cout1237w(0) <= NOT wire_csa_lower_cout;
	loop100 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout1237w1238w1239w(i) <= wire_csa_lower_w_lg_w_lg_cout1237w1238w(i) OR wire_csa_lower_w_lg_cout1236w(i);
	END GENERATE loop100;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(12 DOWNTO 0),
		datab => datab(12 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(25 DOWNTO 13),
		datab => datab(25 DOWNTO 13),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(25 DOWNTO 13),
		datab => datab(25 DOWNTO 13),
		result => wire_csa_upper1_result
	  );

 END RTL; --fplog_altfp_log_csa_p1e

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_add_sub 27 lpm_mult 4 lpm_mux 5 reg 531 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_range_reduction_uqd IS 
	 PORT 
	 ( 
		 a0_in	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 aclr	:	IN  STD_LOGIC := '0';
		 almostlog	:	OUT  STD_LOGIC_VECTOR (38 DOWNTO 0);
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC;
		 y0_in	:	IN  STD_LOGIC_VECTOR (24 DOWNTO 0);
		 z	:	OUT  STD_LOGIC_VECTOR (25 DOWNTO 0)
	 ); 
 END fplog_range_reduction_uqd;

 ARCHITECTURE RTL OF fplog_range_reduction_uqd IS

	 SIGNAL  wire_add0_1_datab	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add0_1_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add0_2_datab	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add0_2_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add0_3_datab	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add0_3_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add1_1_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add1_2_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_add1_3_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_sub1_1_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_sub1_2_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_sub1_3_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL	 A_pipe0_reg0	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 A_pipe0_reg1	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 A_pipe0_reg2	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 A_wire1_reg0	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 A_wire2_reg0	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 A_wire3_reg0	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 B_wire1_reg0	:	STD_LOGIC_VECTOR(20 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 B_wire2_reg0	:	STD_LOGIC_VECTOR(26 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 B_wire3_reg0	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 P_pipe0_reg0	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 P_pipe1_reg0	:	STD_LOGIC_VECTOR(28 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 P_pipe2_reg0	:	STD_LOGIC_VECTOR(28 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 P_pipe3_reg0	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_pipe22_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_pipe23_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_pipe24_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_wire1_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_wire2_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_wire3_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Z_wire1_reg0	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Z_wire2_reg0	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Z_wire3_reg0	:	STD_LOGIC_VECTOR(28 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_mult0_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_mult1_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_mult2_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_mult3_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_InvTable0_data	:	STD_LOGIC_VECTOR (191 DOWNTO 0);
	 SIGNAL  wire_InvTable0_data_2d	:	STD_LOGIC_2D(31 DOWNTO 0, 5 DOWNTO 0);
	 SIGNAL  wire_InvTable0_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_LogTable0_data	:	STD_LOGIC_VECTOR (1247 DOWNTO 0);
	 SIGNAL  wire_LogTable0_data_2d	:	STD_LOGIC_2D(31 DOWNTO 0, 38 DOWNTO 0);
	 SIGNAL  wire_LogTable0_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_LogTable1_data	:	STD_LOGIC_VECTOR (559 DOWNTO 0);
	 SIGNAL  wire_LogTable1_data_2d	:	STD_LOGIC_2D(15 DOWNTO 0, 34 DOWNTO 0);
	 SIGNAL  wire_LogTable1_result	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_LogTable2_data	:	STD_LOGIC_VECTOR (511 DOWNTO 0);
	 SIGNAL  wire_LogTable2_data_2d	:	STD_LOGIC_2D(15 DOWNTO 0, 31 DOWNTO 0);
	 SIGNAL  wire_LogTable2_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_LogTable3_data	:	STD_LOGIC_VECTOR (463 DOWNTO 0);
	 SIGNAL  wire_LogTable3_data_2d	:	STD_LOGIC_2D(15 DOWNTO 0, 28 DOWNTO 0);
	 SIGNAL  wire_LogTable3_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A1_is_not_zero_range999w1017w1018w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_all_zero2_range1089w1093w1097w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_all_zero3_range1166w1170w1174w	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe11_range994w997w998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1078w1079w1080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1082w1083w1084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1086w1087w1088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1155w1156w1157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1159w1160w1161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1163w1164w1165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A1_is_all_zero_range996w1020w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A1_is_not_zero_range999w1016w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A1_is_not_zero_range999w1017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_all_zero2_range1089w1093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_all_zero3_range1166w1170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range994w997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe12_range1074w1075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe12_range1078w1079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe12_range1082w1083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe12_range1086w1087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe13_range1151w1152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe13_range1155w1156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe13_range1159w1160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe13_range1163w1164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w1019w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range984w985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range984w987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range989w990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range989w992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range994w995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  A1_is_all_zero :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A1_is_not_zero :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_all_zero2 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_all_zero3 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_pipe0 :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  A_pipe11 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_pipe12 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_pipe13 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_wire0 :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  A_wire1 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_wire2 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_wire3 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  B_pad_wire1 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  B_pad_wire2 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  B_pad_wire3 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  B_pipe1 :	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  B_pipe2 :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  B_pipe3 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  B_wire1 :	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  B_wire2 :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  B_wire3 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  epsZ_pad_wire1 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  epsZ_pad_wire2 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  epsZ_pad_wire3 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  epsZ_wire1 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  epsZ_wire2 :	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  epsZ_wire3 :	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  InvA0 :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  L_wire0 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  L_wire1 :	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  L_wire2 :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  L_wire3 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  mux0_data0 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  mux0_data1 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  P_pad_wire1 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  P_pad_wire2 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  P_pad_wire3 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  P_pipe0 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  P_pipe1 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  P_pipe2 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  P_pipe3 :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  P_wire0 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  P_wire1 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  P_wire2 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  P_wire3 :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  S_pipe11 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_pipe12 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_pipe13 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_pipe22 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_pipe23 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_pipe24 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_wire1 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_wire2 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_wire3 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_wire4 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  Z_pipe1 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Z_pipe2 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  Z_pipe3 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  Z_wire1 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Z_wire2 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  Z_wire3 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  Z_wire4 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  ZM_wire1 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  ZM_wire2 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  ZM_wire3 :	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_all_zero_range980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_all_zero_range986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_all_zero_range991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_all_zero_range996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_not_zero_range982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_not_zero_range988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_not_zero_range993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_not_zero_range999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero2_range1076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero2_range1081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero2_range1085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero2_range1089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero3_range1153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero3_range1158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero3_range1162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero3_range1166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe11_range984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe11_range989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe11_range994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe12_range1074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe12_range1078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe12_range1082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe12_range1086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe13_range1151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe13_range1155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe13_range1159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe13_range1163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  fplog_altfp_log_csa_s0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(38 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(38 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(38 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_k0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(30 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_r0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(28 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(28 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(28 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_o0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(25 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_l1e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(30 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_s1e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(28 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(28 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(28 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_p1e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(25 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop101 : FOR i IN 0 TO 30 GENERATE 
		wire_range_reduction_w_lg_w_lg_w_A1_is_not_zero_range999w1017w1018w(i) <= wire_range_reduction_w_lg_w_A1_is_not_zero_range999w1017w(0) AND mux0_data0(i);
	END GENERATE loop101;
	loop102 : FOR i IN 0 TO 30 GENERATE 
		wire_range_reduction_w_lg_w_lg_w_A_all_zero2_range1089w1093w1097w(i) <= wire_range_reduction_w_lg_w_A_all_zero2_range1089w1093w(0) AND Z_pipe2(i);
	END GENERATE loop102;
	loop103 : FOR i IN 0 TO 28 GENERATE 
		wire_range_reduction_w_lg_w_lg_w_A_all_zero3_range1166w1170w1174w(i) <= wire_range_reduction_w_lg_w_A_all_zero3_range1166w1170w(0) AND Z_pipe3(i);
	END GENERATE loop103;
	wire_range_reduction_w_lg_w_lg_w_A_pipe11_range994w997w998w(0) <= wire_range_reduction_w_lg_w_A_pipe11_range994w997w(0) AND wire_range_reduction_w_A1_is_not_zero_range993w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1078w1079w1080w(0) <= wire_range_reduction_w_lg_w_A_pipe12_range1078w1079w(0) AND wire_range_reduction_w_A_all_zero2_range1076w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1082w1083w1084w(0) <= wire_range_reduction_w_lg_w_A_pipe12_range1082w1083w(0) AND wire_range_reduction_w_A_all_zero2_range1081w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1086w1087w1088w(0) <= wire_range_reduction_w_lg_w_A_pipe12_range1086w1087w(0) AND wire_range_reduction_w_A_all_zero2_range1085w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1155w1156w1157w(0) <= wire_range_reduction_w_lg_w_A_pipe13_range1155w1156w(0) AND wire_range_reduction_w_A_all_zero3_range1153w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1159w1160w1161w(0) <= wire_range_reduction_w_lg_w_A_pipe13_range1159w1160w(0) AND wire_range_reduction_w_A_all_zero3_range1158w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1163w1164w1165w(0) <= wire_range_reduction_w_lg_w_A_pipe13_range1163w1164w(0) AND wire_range_reduction_w_A_all_zero3_range1162w(0);
	loop104 : FOR i IN 0 TO 30 GENERATE 
		wire_range_reduction_w_lg_w_A1_is_all_zero_range996w1020w(i) <= wire_range_reduction_w_A1_is_all_zero_range996w(0) AND wire_range_reduction_w1019w(i);
	END GENERATE loop104;
	loop105 : FOR i IN 0 TO 30 GENERATE 
		wire_range_reduction_w_lg_w_A1_is_not_zero_range999w1016w(i) <= wire_range_reduction_w_A1_is_not_zero_range999w(0) AND mux0_data1(i);
	END GENERATE loop105;
	wire_range_reduction_w_lg_w_A1_is_not_zero_range999w1017w(0) <= NOT wire_range_reduction_w_A1_is_not_zero_range999w(0);
	wire_range_reduction_w_lg_w_A_all_zero2_range1089w1093w(0) <= NOT wire_range_reduction_w_A_all_zero2_range1089w(0);
	wire_range_reduction_w_lg_w_A_all_zero3_range1166w1170w(0) <= NOT wire_range_reduction_w_A_all_zero3_range1166w(0);
	wire_range_reduction_w_lg_w_A_pipe11_range994w997w(0) <= NOT wire_range_reduction_w_A_pipe11_range994w(0);
	wire_range_reduction_w_lg_w_A_pipe12_range1074w1075w(0) <= NOT wire_range_reduction_w_A_pipe12_range1074w(0);
	wire_range_reduction_w_lg_w_A_pipe12_range1078w1079w(0) <= NOT wire_range_reduction_w_A_pipe12_range1078w(0);
	wire_range_reduction_w_lg_w_A_pipe12_range1082w1083w(0) <= NOT wire_range_reduction_w_A_pipe12_range1082w(0);
	wire_range_reduction_w_lg_w_A_pipe12_range1086w1087w(0) <= NOT wire_range_reduction_w_A_pipe12_range1086w(0);
	wire_range_reduction_w_lg_w_A_pipe13_range1151w1152w(0) <= NOT wire_range_reduction_w_A_pipe13_range1151w(0);
	wire_range_reduction_w_lg_w_A_pipe13_range1155w1156w(0) <= NOT wire_range_reduction_w_A_pipe13_range1155w(0);
	wire_range_reduction_w_lg_w_A_pipe13_range1159w1160w(0) <= NOT wire_range_reduction_w_A_pipe13_range1159w(0);
	wire_range_reduction_w_lg_w_A_pipe13_range1163w1164w(0) <= NOT wire_range_reduction_w_A_pipe13_range1163w(0);
	loop106 : FOR i IN 0 TO 30 GENERATE 
		wire_range_reduction_w1019w(i) <= wire_range_reduction_w_lg_w_lg_w_A1_is_not_zero_range999w1017w1018w(i) OR wire_range_reduction_w_lg_w_A1_is_not_zero_range999w1016w(i);
	END GENERATE loop106;
	wire_range_reduction_w_lg_w_A_pipe11_range984w985w(0) <= wire_range_reduction_w_A_pipe11_range984w(0) OR wire_range_reduction_w_A1_is_all_zero_range980w(0);
	wire_range_reduction_w_lg_w_A_pipe11_range984w987w(0) <= wire_range_reduction_w_A_pipe11_range984w(0) OR wire_range_reduction_w_A1_is_not_zero_range982w(0);
	wire_range_reduction_w_lg_w_A_pipe11_range989w990w(0) <= wire_range_reduction_w_A_pipe11_range989w(0) OR wire_range_reduction_w_A1_is_all_zero_range986w(0);
	wire_range_reduction_w_lg_w_A_pipe11_range989w992w(0) <= wire_range_reduction_w_A_pipe11_range989w(0) OR wire_range_reduction_w_A1_is_not_zero_range988w(0);
	wire_range_reduction_w_lg_w_A_pipe11_range994w995w(0) <= wire_range_reduction_w_A_pipe11_range994w(0) OR wire_range_reduction_w_A1_is_all_zero_range991w(0);
	A1_is_all_zero <= ( wire_range_reduction_w_lg_w_A_pipe11_range994w995w & wire_range_reduction_w_lg_w_A_pipe11_range989w990w & wire_range_reduction_w_lg_w_A_pipe11_range984w985w & A_pipe11(0));
	A1_is_not_zero <= ( wire_range_reduction_w_lg_w_lg_w_A_pipe11_range994w997w998w & wire_range_reduction_w_lg_w_A_pipe11_range989w992w & wire_range_reduction_w_lg_w_A_pipe11_range984w987w & A_pipe11(0));
	A_all_zero2 <= ( wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1086w1087w1088w & wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1082w1083w1084w & wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1078w1079w1080w & wire_range_reduction_w_lg_w_A_pipe12_range1074w1075w);
	A_all_zero3 <= ( wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1163w1164w1165w & wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1159w1160w1161w & wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1155w1156w1157w & wire_range_reduction_w_lg_w_A_pipe13_range1151w1152w);
	A_pipe0 <= a0_in;
	A_pipe11 <= A_wire1_reg0;
	A_pipe12 <= A_wire2_reg0;
	A_pipe13 <= A_wire3_reg0;
	A_wire0 <= A_pipe0_reg2;
	A_wire1 <= Z_wire1(24 DOWNTO 21);
	A_wire2 <= Z_wire2(30 DOWNTO 27);
	A_wire3 <= Z_wire3(28 DOWNTO 25);
	almostlog <= S_wire4;
	B_pad_wire1 <= ( "0" & B_pipe1 & "000000000");
	B_pad_wire2 <= ( "0" & B_pipe2 & "0");
	B_pad_wire3 <= ( "0" & B_pipe3);
	B_pipe1 <= B_wire1_reg0;
	B_pipe2 <= B_wire2_reg0;
	B_pipe3 <= B_wire3_reg0;
	B_wire1 <= Z_wire1(20 DOWNTO 0);
	B_wire2 <= Z_wire2(26 DOWNTO 0);
	B_wire3 <= Z_wire3(24 DOWNTO 0);
	epsZ_pad_wire1 <= epsZ_wire1(30 DOWNTO 0);
	epsZ_pad_wire2 <= epsZ_wire2(39 DOWNTO 11);
	epsZ_pad_wire3 <= epsZ_wire3(40 DOWNTO 15);
	epsZ_wire1 <= wire_range_reduction_w_lg_w_A1_is_all_zero_range996w1020w;
	epsZ_wire2 <= ( "0" & wire_range_reduction_w_lg_w_A_all_zero2_range1089w1093w & "0000000" & wire_range_reduction_w_lg_w_lg_w_A_all_zero2_range1089w1093w1097w);
	epsZ_wire3 <= ( "0" & wire_range_reduction_w_lg_w_A_all_zero3_range1166w1170w & "0000000000" & wire_range_reduction_w_lg_w_lg_w_A_all_zero3_range1166w1170w1174w);
	InvA0 <= wire_InvTable0_result;
	L_wire0 <= wire_LogTable0_result;
	L_wire1 <= wire_LogTable1_result;
	L_wire2 <= wire_LogTable2_result;
	L_wire3 <= wire_LogTable3_result;
	mux0_data0 <= ( "1" & "0000" & Z_pipe1 & "0");
	mux0_data1 <= ( "0" & "1" & "0000" & Z_pipe1);
	P_pad_wire1 <= ( "0" & P_wire1 & "0");
	P_pad_wire2 <= ( "0000" & P_wire2(28 DOWNTO 4));
	P_pad_wire3 <= ( "0000000" & P_wire3(22 DOWNTO 4));
	P_pipe0 <= wire_mult0_result;
	P_pipe1 <= wire_mult1_result;
	P_pipe2 <= wire_mult2_result;
	P_pipe3 <= wire_mult3_result;
	P_wire0 <= P_pipe0_reg0;
	P_wire1 <= P_pipe1_reg0;
	P_wire2 <= P_pipe2_reg0;
	P_wire3 <= P_pipe3_reg0;
	S_pipe11 <= S_wire1_reg0;
	S_pipe12 <= S_wire2_reg0;
	S_pipe13 <= S_wire3_reg0;
	S_pipe22 <= wire_add0_1_result;
	S_pipe23 <= wire_add0_2_result;
	S_pipe24 <= wire_add0_3_result;
	S_wire1 <= L_wire0;
	S_wire2 <= S_pipe22_reg0;
	S_wire3 <= S_pipe23_reg0;
	S_wire4 <= S_pipe24_reg0;
	z <= Z_wire4;
	Z_pipe1 <= Z_wire1_reg0;
	Z_pipe2 <= Z_wire2_reg0;
	Z_pipe3 <= Z_wire3_reg0;
	Z_wire1 <= P_wire0(24 DOWNTO 0);
	Z_wire2 <= wire_sub1_1_result;
	Z_wire3 <= wire_sub1_2_result;
	Z_wire4 <= wire_sub1_3_result;
	ZM_wire1 <= Z_wire1;
	ZM_wire2 <= Z_wire2(30 DOWNTO 6);
	ZM_wire3 <= Z_wire3(28 DOWNTO 10);
	wire_range_reduction_w_A1_is_all_zero_range980w(0) <= A1_is_all_zero(0);
	wire_range_reduction_w_A1_is_all_zero_range986w(0) <= A1_is_all_zero(1);
	wire_range_reduction_w_A1_is_all_zero_range991w(0) <= A1_is_all_zero(2);
	wire_range_reduction_w_A1_is_all_zero_range996w(0) <= A1_is_all_zero(3);
	wire_range_reduction_w_A1_is_not_zero_range982w(0) <= A1_is_not_zero(0);
	wire_range_reduction_w_A1_is_not_zero_range988w(0) <= A1_is_not_zero(1);
	wire_range_reduction_w_A1_is_not_zero_range993w(0) <= A1_is_not_zero(2);
	wire_range_reduction_w_A1_is_not_zero_range999w(0) <= A1_is_not_zero(3);
	wire_range_reduction_w_A_all_zero2_range1076w(0) <= A_all_zero2(0);
	wire_range_reduction_w_A_all_zero2_range1081w(0) <= A_all_zero2(1);
	wire_range_reduction_w_A_all_zero2_range1085w(0) <= A_all_zero2(2);
	wire_range_reduction_w_A_all_zero2_range1089w(0) <= A_all_zero2(3);
	wire_range_reduction_w_A_all_zero3_range1153w(0) <= A_all_zero3(0);
	wire_range_reduction_w_A_all_zero3_range1158w(0) <= A_all_zero3(1);
	wire_range_reduction_w_A_all_zero3_range1162w(0) <= A_all_zero3(2);
	wire_range_reduction_w_A_all_zero3_range1166w(0) <= A_all_zero3(3);
	wire_range_reduction_w_A_pipe11_range984w(0) <= A_pipe11(1);
	wire_range_reduction_w_A_pipe11_range989w(0) <= A_pipe11(2);
	wire_range_reduction_w_A_pipe11_range994w(0) <= A_pipe11(3);
	wire_range_reduction_w_A_pipe12_range1074w(0) <= A_pipe12(0);
	wire_range_reduction_w_A_pipe12_range1078w(0) <= A_pipe12(1);
	wire_range_reduction_w_A_pipe12_range1082w(0) <= A_pipe12(2);
	wire_range_reduction_w_A_pipe12_range1086w(0) <= A_pipe12(3);
	wire_range_reduction_w_A_pipe13_range1151w(0) <= A_pipe13(0);
	wire_range_reduction_w_A_pipe13_range1155w(0) <= A_pipe13(1);
	wire_range_reduction_w_A_pipe13_range1159w(0) <= A_pipe13(2);
	wire_range_reduction_w_A_pipe13_range1163w(0) <= A_pipe13(3);
	wire_add0_1_datab <= ( "0000" & L_wire1);
	add0_1 :  fplog_altfp_log_csa_s0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => S_pipe11,
		datab => wire_add0_1_datab,
		result => wire_add0_1_result
	  );
	wire_add0_2_datab <= ( "0000000" & L_wire2);
	add0_2 :  fplog_altfp_log_csa_s0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => S_pipe12,
		datab => wire_add0_2_datab,
		result => wire_add0_2_result
	  );
	wire_add0_3_datab <= ( "0000000000" & L_wire3);
	add0_3 :  fplog_altfp_log_csa_s0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => S_pipe13,
		datab => wire_add0_3_datab,
		result => wire_add0_3_result
	  );
	add1_1 :  fplog_altfp_log_csa_k0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => B_pad_wire1,
		datab => epsZ_pad_wire1,
		result => wire_add1_1_result
	  );
	add1_2 :  fplog_altfp_log_csa_r0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => B_pad_wire2,
		datab => epsZ_pad_wire2,
		result => wire_add1_2_result
	  );
	add1_3 :  fplog_altfp_log_csa_o0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => B_pad_wire3,
		datab => epsZ_pad_wire3,
		result => wire_add1_3_result
	  );
	sub1_1 :  fplog_altfp_log_csa_l1e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_add1_1_result,
		datab => P_pad_wire1,
		result => wire_sub1_1_result
	  );
	sub1_2 :  fplog_altfp_log_csa_s1e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_add1_2_result,
		datab => P_pad_wire2,
		result => wire_sub1_2_result
	  );
	sub1_3 :  fplog_altfp_log_csa_p1e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_add1_3_result,
		datab => P_pad_wire3,
		result => wire_sub1_3_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_pipe0_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_pipe0_reg0 <= A_pipe0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_pipe0_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_pipe0_reg1 <= A_pipe0_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_pipe0_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_pipe0_reg2 <= A_pipe0_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_wire1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_wire1_reg0 <= A_wire1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_wire2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_wire2_reg0 <= A_wire2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_wire3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_wire3_reg0 <= A_wire3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN B_wire1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN B_wire1_reg0 <= B_wire1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN B_wire2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN B_wire2_reg0 <= B_wire2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN B_wire3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN B_wire3_reg0 <= B_wire3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN P_pipe0_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN P_pipe0_reg0 <= P_pipe0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN P_pipe1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN P_pipe1_reg0 <= P_pipe1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN P_pipe2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN P_pipe2_reg0 <= P_pipe2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN P_pipe3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN P_pipe3_reg0 <= P_pipe3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_pipe22_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_pipe22_reg0 <= S_pipe22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_pipe23_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_pipe23_reg0 <= S_pipe23;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_pipe24_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_pipe24_reg0 <= S_pipe24;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_wire1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_wire1_reg0 <= S_wire1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_wire2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_wire2_reg0 <= S_wire2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_wire3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_wire3_reg0 <= S_wire3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Z_wire1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Z_wire1_reg0 <= Z_wire1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Z_wire2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Z_wire2_reg0 <= Z_wire2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Z_wire3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Z_wire3_reg0 <= Z_wire3;
			END IF;
		END IF;
	END PROCESS;
	mult0 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 6,
		LPM_WIDTHB => 25,
		LPM_WIDTHP => 31
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => InvA0,
		datab => y0_in,
		result => wire_mult0_result
	  );
	mult1 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 4,
		LPM_WIDTHB => 25,
		LPM_WIDTHP => 29
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => A_wire1,
		datab => ZM_wire1,
		result => wire_mult1_result
	  );
	mult2 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 4,
		LPM_WIDTHB => 25,
		LPM_WIDTHP => 29
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => A_wire2,
		datab => ZM_wire2,
		result => wire_mult2_result
	  );
	mult3 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 4,
		LPM_WIDTHB => 19,
		LPM_WIDTHP => 23
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => A_wire3,
		datab => ZM_wire3,
		result => wire_mult3_result
	  );
	wire_InvTable0_data <= ( "100001" & "100010" & "100010" & "100011" & "100011" & "100100" & "100100" & "100101" & "100110" & "100110" & "100111" & "101000" & "101001" & "101001" & "101010" & "101011" & "010110" & "010111" & "010111" & "011000" & "011000" & "011001" & "011001" & "011010" & "011011" & "011011" & "011100" & "011101" & "011110" & "011111" & "100000" & "100000");
	loop107 : FOR i IN 0 TO 31 GENERATE
		loop108 : FOR j IN 0 TO 5 GENERATE
			wire_InvTable0_data_2d(i, j) <= wire_InvTable0_data(i*6+j);
		END GENERATE loop108;
	END GENERATE loop107;
	InvTable0 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 32,
		LPM_WIDTH => 6,
		LPM_WIDTHS => 5
	  )
	  PORT MAP ( 
		data => wire_InvTable0_data_2d,
		result => wire_InvTable0_result,
		sel => a0_in
	  );
	wire_LogTable0_data <= ( "111110000001111101011001001111000110001" & "111100000111101011100111100111111111100" & "111100000111101011100111100111111111100" & "111010010000111100101101011101010001110" & "111010010000111100101101011101010001110" & "111000011101100011111000100100011101011" & "111000011101100011111000100100011101011" & "110110101101010101011010000011111100001" & "110101000000000110011111000111101011001" & "110101000000000110011111000111101011001" & "110011010101101101001010110001100001100" & "110001101110000000010000011100001100110" & "110000001000110111001111001001010100010" & "110000001000110111001111001001010100010" & "101110100110001010001101010100010101001" & "101101000101110001110101000101000111110" & "010111111110101111101000111011110110000" & "010101001000101010111000000111001110001" & "010101001000101010111000000111001110001" & "010010011010010110001000010001001101001" & "010010011010010110001000010001001101001" & "001111110011001000111000110110010110011" & "001111110011001000111000110110010110011" & "001101010010011111011010011110010001010" & "001010110111111010000000110101101010100" & "001010110111111010000000110101101010100" & "001000100010111100011101000001000100111" & "000110010011001101011110010111010101100" & "000100001000010110011000101101011001111" & "000010000010000010101110110001001111001" & "000000000000000000000000000000000000000" & "000000000000000000000000000000000000000");
	loop109 : FOR i IN 0 TO 31 GENERATE
		loop110 : FOR j IN 0 TO 38 GENERATE
			wire_LogTable0_data_2d(i, j) <= wire_LogTable0_data(i*39+j);
		END GENERATE loop110;
	END GENERATE loop109;
	LogTable0 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 32,
		LPM_WIDTH => 39,
		LPM_WIDTHS => 5
	  )
	  PORT MAP ( 
		data => wire_LogTable0_data_2d,
		result => wire_LogTable0_result,
		sel => A_wire0
	  );
	wire_LogTable1_data <= ( "11100110010110111001111001101110111" & "11010101011101111001011010000111110" & "11000100101001010101000010100100111" & "10110011111001001010011110010110101" & "10100011001101010111011010100001011" & "10010010100101111001100101111100011" & "10000010000010101110110001001111001" & "01110001100011110100101110110000010" & "01101001010101111101010100100011000" & "01011000111101011000010111100001101" & "01001000101000111110110001111111101" & "00111000011000101110011100001001100" & "00101000001100100101001111110010110" & "00011000000100100001001000010100010" & "00001000000000100000000010101010111" & "00000000000000000000000000000000000");
	loop111 : FOR i IN 0 TO 15 GENERATE
		loop112 : FOR j IN 0 TO 34 GENERATE
			wire_LogTable1_data_2d(i, j) <= wire_LogTable1_data(i*35+j);
		END GENERATE loop112;
	END GENERATE loop111;
	LogTable1 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 16,
		LPM_WIDTH => 35,
		LPM_WIDTHS => 4
	  )
	  PORT MAP ( 
		data => wire_LogTable1_data_2d,
		result => wire_LogTable1_result,
		sel => A_pipe11
	  );
	wire_LogTable2_data <= ( "11101000110100110011111101101000" & "11011000101101110000111000001100" & "11001000100111001110001110000010" & "10111000100001001011111101000110" & "10101000011011101010000011010111" & "10011000010110101000011110110010" & "10001000010010000111001101010110" & "01111000001110000110001101000000" & "01101000001010100101011011110000" & "01011000000111100100110111100100" & "01001000000101000100011110011011" & "00111000000011000100001110010011" & "00101000000001100100000101001101" & "00011000000000100100000001001000" & "00001000000000000100000000000010" & "00000000000000000000000000000000");
	loop113 : FOR i IN 0 TO 15 GENERATE
		loop114 : FOR j IN 0 TO 31 GENERATE
			wire_LogTable2_data_2d(i, j) <= wire_LogTable2_data(i*32+j);
		END GENERATE loop114;
	END GENERATE loop113;
	LogTable2 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 16,
		LPM_WIDTH => 32,
		LPM_WIDTHS => 4
	  )
	  PORT MAP ( 
		data => wire_LogTable2_data_2d,
		result => wire_LogTable2_result,
		sel => A_pipe12
	  );
	wire_LogTable3_data <= ( "11101000000110100100101111111" & "11011000000101101100101100110" & "11001000000100111000101010001" & "10111000000100001000100111111" & "10101000000011011100100110000" & "10011000000010110100100100011" & "10001000000010010000100011001" & "01111000000001110000100010001" & "01101000000001010100100001011" & "01011000000000111100100000110" & "01001000000000101000100000011" & "00111000000000011000100000001" & "00101000000000001100100000000" & "00011000000000000100100000000" & "00001000000000000000100000000" & "00000000000000000000000000000");
	loop115 : FOR i IN 0 TO 15 GENERATE
		loop116 : FOR j IN 0 TO 28 GENERATE
			wire_LogTable3_data_2d(i, j) <= wire_LogTable3_data(i*29+j);
		END GENERATE loop116;
	END GENERATE loop115;
	LogTable3 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 16,
		LPM_WIDTH => 29,
		LPM_WIDTHS => 4
	  )
	  PORT MAP ( 
		data => wire_LogTable3_data_2d,
		result => wire_LogTable3_result,
		sel => A_pipe13
	  );

 END RTL; --fplog_range_reduction_uqd


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" PIPELINE=1 WIDTH=64 WIDTHAD=6 aclr clk_en clock data q
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" PIPELINE=0 WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END fplog_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --fplog_altpriority_encoder_3v7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END fplog_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --fplog_altpriority_encoder_3e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END fplog_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_w_lg_zero1280w1281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_zero1282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_zero1280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_w_lg_zero1282w1283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_zero	:	STD_LOGIC;
	 COMPONENT  fplog_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder15_w_lg_zero1280w & wire_altpriority_encoder15_w_lg_w_lg_zero1282w1283w);
	altpriority_encoder14 :  fplog_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder14_q
	  );
	wire_altpriority_encoder15_w_lg_w_lg_zero1280w1281w(0) <= wire_altpriority_encoder15_w_lg_zero1280w(0) AND wire_altpriority_encoder15_q(0);
	wire_altpriority_encoder15_w_lg_zero1282w(0) <= wire_altpriority_encoder15_zero AND wire_altpriority_encoder14_q(0);
	wire_altpriority_encoder15_w_lg_zero1280w(0) <= NOT wire_altpriority_encoder15_zero;
	wire_altpriority_encoder15_w_lg_w_lg_zero1282w1283w(0) <= wire_altpriority_encoder15_w_lg_zero1282w(0) OR wire_altpriority_encoder15_w_lg_w_lg_zero1280w1281w(0);
	altpriority_encoder15 :  fplog_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder15_q,
		zero => wire_altpriority_encoder15_zero
	  );

 END RTL; --fplog_altpriority_encoder_6v7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END fplog_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder16_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder17_w_lg_w_lg_zero1298w1299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_w_lg_zero1300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_w_lg_zero1298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_w_lg_w_lg_zero1300w1301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_zero	:	STD_LOGIC;
	 COMPONENT  fplog_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder17_w_lg_zero1298w & wire_altpriority_encoder17_w_lg_w_lg_zero1300w1301w);
	zero <= (wire_altpriority_encoder16_zero AND wire_altpriority_encoder17_zero);
	altpriority_encoder16 :  fplog_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder16_q,
		zero => wire_altpriority_encoder16_zero
	  );
	wire_altpriority_encoder17_w_lg_w_lg_zero1298w1299w(0) <= wire_altpriority_encoder17_w_lg_zero1298w(0) AND wire_altpriority_encoder17_q(0);
	wire_altpriority_encoder17_w_lg_zero1300w(0) <= wire_altpriority_encoder17_zero AND wire_altpriority_encoder16_q(0);
	wire_altpriority_encoder17_w_lg_zero1298w(0) <= NOT wire_altpriority_encoder17_zero;
	wire_altpriority_encoder17_w_lg_w_lg_zero1300w1301w(0) <= wire_altpriority_encoder17_w_lg_zero1300w(0) OR wire_altpriority_encoder17_w_lg_w_lg_zero1298w1299w(0);
	altpriority_encoder17 :  fplog_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder17_q,
		zero => wire_altpriority_encoder17_zero
	  );

 END RTL; --fplog_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END fplog_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_w_lg_zero1271w1272w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_zero1273w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_zero1271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_w_lg_zero1273w1274w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 COMPONENT  fplog_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder13_w_lg_zero1271w & wire_altpriority_encoder13_w_lg_w_lg_zero1273w1274w);
	altpriority_encoder12 :  fplog_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder12_q
	  );
	loop117 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder13_w_lg_w_lg_zero1271w1272w(i) <= wire_altpriority_encoder13_w_lg_zero1271w(0) AND wire_altpriority_encoder13_q(i);
	END GENERATE loop117;
	loop118 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder13_w_lg_zero1273w(i) <= wire_altpriority_encoder13_zero AND wire_altpriority_encoder12_q(i);
	END GENERATE loop118;
	wire_altpriority_encoder13_w_lg_zero1271w(0) <= NOT wire_altpriority_encoder13_zero;
	loop119 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder13_w_lg_w_lg_zero1273w1274w(i) <= wire_altpriority_encoder13_w_lg_zero1273w(i) OR wire_altpriority_encoder13_w_lg_w_lg_zero1271w1272w(i);
	END GENERATE loop119;
	altpriority_encoder13 :  fplog_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );

 END RTL; --fplog_altpriority_encoder_bv7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END fplog_altpriority_encoder_be8;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder18_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder19_w_lg_w_lg_zero1308w1309w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_w_lg_zero1310w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_w_lg_zero1308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_w_lg_w_lg_zero1310w1311w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_zero	:	STD_LOGIC;
	 COMPONENT  fplog_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder19_w_lg_zero1308w & wire_altpriority_encoder19_w_lg_w_lg_zero1310w1311w);
	zero <= (wire_altpriority_encoder18_zero AND wire_altpriority_encoder19_zero);
	altpriority_encoder18 :  fplog_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder18_q,
		zero => wire_altpriority_encoder18_zero
	  );
	loop120 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder19_w_lg_w_lg_zero1308w1309w(i) <= wire_altpriority_encoder19_w_lg_zero1308w(0) AND wire_altpriority_encoder19_q(i);
	END GENERATE loop120;
	loop121 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder19_w_lg_zero1310w(i) <= wire_altpriority_encoder19_zero AND wire_altpriority_encoder18_q(i);
	END GENERATE loop121;
	wire_altpriority_encoder19_w_lg_zero1308w(0) <= NOT wire_altpriority_encoder19_zero;
	loop122 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder19_w_lg_w_lg_zero1310w1311w(i) <= wire_altpriority_encoder19_w_lg_zero1310w(i) OR wire_altpriority_encoder19_w_lg_w_lg_zero1308w1309w(i);
	END GENERATE loop122;
	altpriority_encoder19 :  fplog_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder19_q,
		zero => wire_altpriority_encoder19_zero
	  );

 END RTL; --fplog_altpriority_encoder_be8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_r08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END fplog_altpriority_encoder_r08;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_r08 IS

	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_w_lg_zero1262w1263w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_zero1264w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_zero1262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_w_lg_zero1264w1265w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 COMPONENT  fplog_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder11_w_lg_zero1262w & wire_altpriority_encoder11_w_lg_w_lg_zero1264w1265w);
	altpriority_encoder10 :  fplog_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder10_q
	  );
	loop123 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder11_w_lg_w_lg_zero1262w1263w(i) <= wire_altpriority_encoder11_w_lg_zero1262w(0) AND wire_altpriority_encoder11_q(i);
	END GENERATE loop123;
	loop124 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder11_w_lg_zero1264w(i) <= wire_altpriority_encoder11_zero AND wire_altpriority_encoder10_q(i);
	END GENERATE loop124;
	wire_altpriority_encoder11_w_lg_zero1262w(0) <= NOT wire_altpriority_encoder11_zero;
	loop125 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder11_w_lg_w_lg_zero1264w1265w(i) <= wire_altpriority_encoder11_w_lg_zero1264w(i) OR wire_altpriority_encoder11_w_lg_w_lg_zero1262w1263w(i);
	END GENERATE loop125;
	altpriority_encoder11 :  fplog_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );

 END RTL; --fplog_altpriority_encoder_r08


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_rf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END fplog_altpriority_encoder_rf8;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_rf8 IS

	 SIGNAL  wire_altpriority_encoder20_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder21_w_lg_w_lg_zero1318w1319w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_w_lg_zero1320w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_w_lg_zero1318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_w_lg_w_lg_zero1320w1321w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_zero	:	STD_LOGIC;
	 COMPONENT  fplog_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder21_w_lg_zero1318w & wire_altpriority_encoder21_w_lg_w_lg_zero1320w1321w);
	zero <= (wire_altpriority_encoder20_zero AND wire_altpriority_encoder21_zero);
	altpriority_encoder20 :  fplog_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder20_q,
		zero => wire_altpriority_encoder20_zero
	  );
	loop126 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder21_w_lg_w_lg_zero1318w1319w(i) <= wire_altpriority_encoder21_w_lg_zero1318w(0) AND wire_altpriority_encoder21_q(i);
	END GENERATE loop126;
	loop127 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder21_w_lg_zero1320w(i) <= wire_altpriority_encoder21_zero AND wire_altpriority_encoder20_q(i);
	END GENERATE loop127;
	wire_altpriority_encoder21_w_lg_zero1318w(0) <= NOT wire_altpriority_encoder21_zero;
	loop128 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder21_w_lg_w_lg_zero1320w1321w(i) <= wire_altpriority_encoder21_w_lg_zero1320w(i) OR wire_altpriority_encoder21_w_lg_w_lg_zero1318w1319w(i);
	END GENERATE loop128;
	altpriority_encoder21 :  fplog_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder21_q,
		zero => wire_altpriority_encoder21_zero
	  );

 END RTL; --fplog_altpriority_encoder_rf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_tv8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END fplog_altpriority_encoder_tv8;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_tv8 IS

	 SIGNAL  wire_altpriority_encoder8_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_w_lg_zero1253w1254w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_zero1255w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_zero1253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_w_lg_zero1255w1256w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_zero	:	STD_LOGIC;
	 COMPONENT  fplog_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder9_w_lg_zero1253w & wire_altpriority_encoder9_w_lg_w_lg_zero1255w1256w);
	altpriority_encoder8 :  fplog_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder8_q
	  );
	loop129 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder9_w_lg_w_lg_zero1253w1254w(i) <= wire_altpriority_encoder9_w_lg_zero1253w(0) AND wire_altpriority_encoder9_q(i);
	END GENERATE loop129;
	loop130 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder9_w_lg_zero1255w(i) <= wire_altpriority_encoder9_zero AND wire_altpriority_encoder8_q(i);
	END GENERATE loop130;
	wire_altpriority_encoder9_w_lg_zero1253w(0) <= NOT wire_altpriority_encoder9_zero;
	loop131 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder9_w_lg_w_lg_zero1255w1256w(i) <= wire_altpriority_encoder9_w_lg_zero1255w(i) OR wire_altpriority_encoder9_w_lg_w_lg_zero1253w1254w(i);
	END GENERATE loop131;
	altpriority_encoder9 :  fplog_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder9_q,
		zero => wire_altpriority_encoder9_zero
	  );

 END RTL; --fplog_altpriority_encoder_tv8


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" PIPELINE=0 WIDTH=32 WIDTHAD=5 data q zero
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_te9 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END fplog_altpriority_encoder_te9;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_te9 IS

	 SIGNAL  wire_altpriority_encoder22_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder23_w_lg_w_lg_zero1328w1329w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_w_lg_zero1330w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_w_lg_zero1328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_w_lg_w_lg_zero1330w1331w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_zero	:	STD_LOGIC;
	 COMPONENT  fplog_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder23_w_lg_zero1328w & wire_altpriority_encoder23_w_lg_w_lg_zero1330w1331w);
	zero <= (wire_altpriority_encoder22_zero AND wire_altpriority_encoder23_zero);
	altpriority_encoder22 :  fplog_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder22_q,
		zero => wire_altpriority_encoder22_zero
	  );
	loop132 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder23_w_lg_w_lg_zero1328w1329w(i) <= wire_altpriority_encoder23_w_lg_zero1328w(0) AND wire_altpriority_encoder23_q(i);
	END GENERATE loop132;
	loop133 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder23_w_lg_zero1330w(i) <= wire_altpriority_encoder23_zero AND wire_altpriority_encoder22_q(i);
	END GENERATE loop133;
	wire_altpriority_encoder23_w_lg_zero1328w(0) <= NOT wire_altpriority_encoder23_zero;
	loop134 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder23_w_lg_w_lg_zero1330w1331w(i) <= wire_altpriority_encoder23_w_lg_zero1330w(i) OR wire_altpriority_encoder23_w_lg_w_lg_zero1328w1329w(i);
	END GENERATE loop134;
	altpriority_encoder23 :  fplog_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder23_q,
		zero => wire_altpriority_encoder23_zero
	  );

 END RTL; --fplog_altpriority_encoder_te9

--synthesis_resources = reg 6 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_uja IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0)
	 ); 
 END fplog_altpriority_encoder_uja;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_uja IS

	 SIGNAL  wire_altpriority_encoder6_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_w_lg_zero1243w1244w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_zero1245w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_zero1243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_w_lg_zero1245w1246w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_zero	:	STD_LOGIC;
	 SIGNAL	 pipeline_q_dffe	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  tmp_q_wire :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 COMPONENT  fplog_altpriority_encoder_tv8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altpriority_encoder_te9
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= pipeline_q_dffe;
	tmp_q_wire <= ( wire_altpriority_encoder7_w_lg_zero1243w & wire_altpriority_encoder7_w_lg_w_lg_zero1245w1246w);
	altpriority_encoder6 :  fplog_altpriority_encoder_tv8
	  PORT MAP ( 
		data => data(31 DOWNTO 0),
		q => wire_altpriority_encoder6_q
	  );
	loop135 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder7_w_lg_w_lg_zero1243w1244w(i) <= wire_altpriority_encoder7_w_lg_zero1243w(0) AND wire_altpriority_encoder7_q(i);
	END GENERATE loop135;
	loop136 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder7_w_lg_zero1245w(i) <= wire_altpriority_encoder7_zero AND wire_altpriority_encoder6_q(i);
	END GENERATE loop136;
	wire_altpriority_encoder7_w_lg_zero1243w(0) <= NOT wire_altpriority_encoder7_zero;
	loop137 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder7_w_lg_w_lg_zero1245w1246w(i) <= wire_altpriority_encoder7_w_lg_zero1245w(i) OR wire_altpriority_encoder7_w_lg_w_lg_zero1243w1244w(i);
	END GENERATE loop137;
	altpriority_encoder7 :  fplog_altpriority_encoder_te9
	  PORT MAP ( 
		data => data(63 DOWNTO 32),
		q => wire_altpriority_encoder7_q,
		zero => wire_altpriority_encoder7_zero
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN pipeline_q_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN pipeline_q_dffe <= tmp_q_wire;
			END IF;
		END IF;
	END PROCESS;

 END RTL; --fplog_altpriority_encoder_uja


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 16.1 cbx_altpriority_encoder 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altpriority_encoder_q08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END fplog_altpriority_encoder_q08;

 ARCHITECTURE RTL OF fplog_altpriority_encoder_q08 IS

	 SIGNAL  wire_altpriority_encoder24_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_w_lg_w_lg_zero1338w1339w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_w_lg_zero1340w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_w_lg_zero1338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_w_lg_w_lg_zero1340w1341w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_zero	:	STD_LOGIC;
	 COMPONENT  fplog_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder25_w_lg_zero1338w & wire_altpriority_encoder25_w_lg_w_lg_zero1340w1341w);
	altpriority_encoder24 :  fplog_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder24_q
	  );
	loop138 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder25_w_lg_w_lg_zero1338w1339w(i) <= wire_altpriority_encoder25_w_lg_zero1338w(0) AND wire_altpriority_encoder25_q(i);
	END GENERATE loop138;
	loop139 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder25_w_lg_zero1340w(i) <= wire_altpriority_encoder25_zero AND wire_altpriority_encoder24_q(i);
	END GENERATE loop139;
	wire_altpriority_encoder25_w_lg_zero1338w(0) <= NOT wire_altpriority_encoder25_zero;
	loop140 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder25_w_lg_w_lg_zero1340w1341w(i) <= wire_altpriority_encoder25_w_lg_zero1340w(i) OR wire_altpriority_encoder25_w_lg_w_lg_zero1338w1339w(i);
	END GENERATE loop140;
	altpriority_encoder25 :  fplog_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder25_q,
		zero => wire_altpriority_encoder25_zero
	  );

 END RTL; --fplog_altpriority_encoder_q08

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = altsquare 1 lpm_add_sub 42 lpm_mult 5 lpm_mux 5 mux21 31 reg 1563 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fplog_altfp_log_n6b IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 nan	:	OUT  STD_LOGIC;
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END fplog_altfp_log_n6b;

 ARCHITECTURE RTL OF fplog_altfp_log_n6b IS

	 SIGNAL  wire_Lshiftsmall_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_data	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_distance	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_E_w_lg_q189w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_result	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_exp_nan_result	:	STD_LOGIC;
	 SIGNAL  wire_exp_zero_result	:	STD_LOGIC;
	 SIGNAL  wire_man_inf_result	:	STD_LOGIC;
	 SIGNAL  wire_man_nan_result	:	STD_LOGIC;
	 SIGNAL  wire_add1_dataa	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add1_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add2_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add2_datab	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add2_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_exp_biase_sub_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub1_dataa	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_sub1_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_sub2_dataa	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub2_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub3_dataa	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_sub3_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_sub3_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_sub4_datab	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_sub4_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_sub5_dataa	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub5_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub5_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub6_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub6_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_range_reduction_almostlog	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_range_reduction_z	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_E_data	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_E_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_lzoc_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_lzoc_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_squarer_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL	 absELog2_pipe_reg0	:	STD_LOGIC_VECTOR(34 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absELog2_pipe_reg1	:	STD_LOGIC_VECTOR(34 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absELog2_pipe_reg2	:	STD_LOGIC_VECTOR(34 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg0	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg1	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg2	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg3	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg4	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg5	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg6	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg7	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg8	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg9	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0s_pipe1_reg0	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0s_pipe1_reg1	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0s_pipe1_reg2	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0s_pipe1_reg3	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0s_reg0	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 almostLog_pipe_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 almostLog_pipe_reg1	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 almostLog_pipe_reg2	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 doRR_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 doRR_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg0	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg1	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg4	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg5	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg6	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg7	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg8	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg9	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E_normal_pipe_reg0	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_is_ebiase_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_is_ebiase_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_is_ebiase_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg10	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg11	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg12	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg13	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg14	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg15	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg16	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg17	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg10	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg11	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg12	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg13	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg14	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg15	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg16	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg17	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg10	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg11	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg12	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg13	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg14	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg15	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg16	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg17	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg10	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg11	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg12	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg13	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg14	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg15	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg16	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg17	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Log_normal_normd_pipe_reg0	:	STD_LOGIC_VECTOR(46 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Log_normal_reg0	:	STD_LOGIC_VECTOR(46 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Log_small_normd_pipe_reg0	:	STD_LOGIC_VECTOR(26 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Log_small_normd_pipe_reg1	:	STD_LOGIC_VECTOR(26 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Lshiftval_reg0	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Lshiftval_reg1	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Lshiftval_reg2	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Lshiftval_reg3	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg0	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg1	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg2	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg3	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg4	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg5	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg6	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg7	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg8	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg9	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg0	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg1	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg2	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg3	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg4	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg5	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg6	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg7	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_data_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_data_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_data_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe3_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe3_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe3_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe3_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe3_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Z2o2_pipe_reg0	:	STD_LOGIC_VECTOR(13 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Z2o2_small_s_pipe_reg0	:	STD_LOGIC_VECTOR(13 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Zfinal_reg0	:	STD_LOGIC_VECTOR(25 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Zfinal_reg1	:	STD_LOGIC_VECTOR(25 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_addsub1_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_addsub2_add_sub	:	STD_LOGIC;
	 SIGNAL  wire_addsub2_result	:	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  wire_mult1_result	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL	wire_mux_result0a_dataout	:	STD_LOGIC_VECTOR(30 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_doRR_pipe125w126w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_First_bit9w83w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_small_flag206w215w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_small_flag206w207w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sR_pipe188w89w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sR_pipe292w93w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range42w43w44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range46w47w48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range50w51w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range54w55w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range58w59w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range62w63w64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range66w67w68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_exp_data_range31w33w34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_Log_small_range149w154w194w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_Log_small_range150w198w199w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_sR254w255w256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_doRR_pipe124w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_lg_First_bit82w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_w_lg_small_flag214w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_small_flag204w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR_pipe187w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR_pipe291w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range13w15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range16w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range19w21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range22w24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range25w27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range28w30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_g_range228w229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range149w192w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range150w197w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_doRR111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_doRR_pipe125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_E_normal212w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_all_zero240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_First_bit9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_is_one247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_all_zero241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_small_flag206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR_pipe188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR_pipe292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR_pipe3179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range38w39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range42w43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range46w47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range50w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range54w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range58w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range62w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range66w67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range31w33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range149w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range150w198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_input_is_one247w248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_input_is_zero244w245w246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_input_is_zero244w245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sR254w255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_is_zero244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_g_range220w221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_g_range223w224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_g_range226w227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range150w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range150w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_First_bit96w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  absE :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  absELog2 :	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  absELog2_pad :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  absELog2_pipe :	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  absZ0 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  absZ0_pipe :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  absZ0s :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  absZ0s_pipe1 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  absZ0s_pipe2 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  almostLog :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  almostLog_pipe :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  data_exp_is_ebiase :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  doRR :	STD_LOGIC;
	 SIGNAL  doRR_pipe :	STD_LOGIC;
	 SIGNAL  E0 :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  E0_is_zero :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  E0_pipe :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  E0_sub :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  E0offset :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  E_normal :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  E_normal_pipe :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  E_small :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  EFR :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  ER :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_all_one :	STD_LOGIC;
	 SIGNAL  exp_all_zero :	STD_LOGIC;
	 SIGNAL  exp_biase :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_data :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_is_ebiase :	STD_LOGIC;
	 SIGNAL  exp_is_ebiase_pipe :	STD_LOGIC;
	 SIGNAL  First_bit :	STD_LOGIC;
	 SIGNAL  input_is_infinity :	STD_LOGIC;
	 SIGNAL  input_is_infinity_pipe :	STD_LOGIC;
	 SIGNAL  input_is_nan :	STD_LOGIC;
	 SIGNAL  input_is_nan_pipe :	STD_LOGIC;
	 SIGNAL  input_is_one :	STD_LOGIC;
	 SIGNAL  input_is_one_pipe :	STD_LOGIC;
	 SIGNAL  input_is_zero :	STD_LOGIC;
	 SIGNAL  input_is_zero_pipe :	STD_LOGIC;
	 SIGNAL  Log1p_normal :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  Log2 :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Log_g :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Log_normal :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  Log_normal_normd :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  Log_normal_normd_pipe :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  Log_normal_pipe :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  Log_small :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  Log_small1 :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Log_small2 :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Log_small_normd :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Log_small_normd_pipe :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  LogF_normal :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  LogF_normal_pad :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  Lshiftval :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  lzo :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  lzo_pipe1 :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  lzo_pipe2 :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  man_above_half :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  man_all_zero :	STD_LOGIC;
	 SIGNAL  man_below_half :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  man_data :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_not_zero :	STD_LOGIC;
	 SIGNAL  pfinal_s :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  round :	STD_LOGIC;
	 SIGNAL  Rshiftval :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sign_data :	STD_LOGIC;
	 SIGNAL  sign_data_pipe :	STD_LOGIC;
	 SIGNAL  small_flag :	STD_LOGIC;
	 SIGNAL  small_flag_pipe :	STD_LOGIC;
	 SIGNAL  squarerIn :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  squarerIn0 :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  squarerIn1 :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  sR :	STD_LOGIC;
	 SIGNAL  sR_pipe1 :	STD_LOGIC;
	 SIGNAL  sR_pipe2 :	STD_LOGIC;
	 SIGNAL  sR_pipe3 :	STD_LOGIC;
	 SIGNAL  sticky :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w203w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Y0 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Z2o2 :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  Z2o2_pipe :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  Z2o2_small :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  Z2o2_small_s :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  Z2o2_small_s_pipe :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  Z_small :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  Zfinal :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  Zfinal_pipe :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_g_range220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_g_range223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_g_range228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_g_range226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_normal_normd_range205w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_Log_small_range193w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_Log_small_range191w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_Log_small_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_small_range196w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_Log_small_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_range222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_range225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Y0_range86w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_Y0_range95w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 COMPONENT  fplog_altbarrel_shift_itd
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altbarrel_shift_qab
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(63 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altbarrel_shift_51e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_and_or_h9b
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_and_or_v6b
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_and_or_c8b
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(22 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_s0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(38 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(38 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(38 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_k0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(30 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_0nc
	 PORT
	 ( 
		dataa	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_d4b
	 PORT
	 ( 
		dataa	:	IN  STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(11 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_umc
	 PORT
	 ( 
		dataa	:	IN  STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_nlf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(25 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altfp_log_csa_8kf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_range_reduction_uqd
	 PORT
	 ( 
		a0_in	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		aclr	:	IN  STD_LOGIC := '0';
		almostlog	:	OUT  STD_LOGIC_VECTOR(38 DOWNTO 0);
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC;
		y0_in	:	IN  STD_LOGIC_VECTOR(24 DOWNTO 0);
		z	:	OUT  STD_LOGIC_VECTOR(25 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altpriority_encoder_uja
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  fplog_altpriority_encoder_q08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altsquare
	 GENERIC 
	 (
		DATA_WIDTH	:	NATURAL;
		PIPELINE	:	NATURAL;
		REPRESENTATION	:	STRING := "UNSIGNED";
		RESULT_ALIGNMENT	:	STRING := "LSB";
		RESULT_WIDTH	:	NATURAL;
		lpm_type	:	STRING := "altsquare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clock	:	IN STD_LOGIC := '1';
		data	:	IN STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
		ena	:	IN STD_LOGIC := '1';
		result	:	OUT STD_LOGIC_VECTOR(RESULT_WIDTH-1 DOWNTO 0)
		-- sclr	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop141 : FOR i IN 0 TO 12 GENERATE 
		wire_w_lg_w_lg_doRR_pipe125w126w(i) <= wire_w_lg_doRR_pipe125w(0) AND squarerIn0(i);
	END GENERATE loop141;
	loop142 : FOR i IN 0 TO 24 GENERATE 
		wire_w_lg_w_lg_First_bit9w83w(i) <= wire_w_lg_First_bit9w(0) AND man_below_half(i);
	END GENERATE loop142;
	loop143 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_small_flag206w215w(i) <= wire_w_lg_small_flag206w(0) AND wire_sub6_result(i);
	END GENERATE loop143;
	loop144 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_w_lg_small_flag206w207w(i) <= wire_w_lg_small_flag206w(0) AND wire_w_Log_normal_normd_range205w(i);
	END GENERATE loop144;
	loop145 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_w_lg_sR_pipe188w89w(i) <= wire_w_lg_sR_pipe188w(0) AND wire_w_Y0_range86w(i);
	END GENERATE loop145;
	loop146 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_sR_pipe292w93w(i) <= wire_w_lg_sR_pipe292w(0) AND E0(i);
	END GENERATE loop146;
	wire_w_lg_w_lg_w_E0_range42w43w44w(0) <= wire_w_lg_w_E0_range42w43w(0) AND wire_w_E0_is_zero_range40w(0);
	wire_w_lg_w_lg_w_E0_range46w47w48w(0) <= wire_w_lg_w_E0_range46w47w(0) AND wire_w_E0_is_zero_range45w(0);
	wire_w_lg_w_lg_w_E0_range50w51w52w(0) <= wire_w_lg_w_E0_range50w51w(0) AND wire_w_E0_is_zero_range49w(0);
	wire_w_lg_w_lg_w_E0_range54w55w56w(0) <= wire_w_lg_w_E0_range54w55w(0) AND wire_w_E0_is_zero_range53w(0);
	wire_w_lg_w_lg_w_E0_range58w59w60w(0) <= wire_w_lg_w_E0_range58w59w(0) AND wire_w_E0_is_zero_range57w(0);
	wire_w_lg_w_lg_w_E0_range62w63w64w(0) <= wire_w_lg_w_E0_range62w63w(0) AND wire_w_E0_is_zero_range61w(0);
	wire_w_lg_w_lg_w_E0_range66w67w68w(0) <= wire_w_lg_w_E0_range66w67w(0) AND wire_w_E0_is_zero_range65w(0);
	wire_w_lg_w_lg_w_exp_data_range31w33w34w(0) <= wire_w_lg_w_exp_data_range31w33w(0) AND wire_w_data_exp_is_ebiase_range29w(0);
	loop147 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_w_lg_w_Log_small_range149w154w194w(i) <= wire_w_lg_w_Log_small_range149w154w(0) AND wire_w_Log_small_range193w(i);
	END GENERATE loop147;
	loop148 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_w_lg_w_Log_small_range150w198w199w(i) <= wire_w_lg_w_Log_small_range150w198w(0) AND Log_small1(i);
	END GENERATE loop148;
	wire_w_lg_w_lg_w_lg_sR254w255w256w(0) <= wire_w_lg_w_lg_sR254w255w(0) AND wire_w_lg_input_is_one247w(0);
	loop149 : FOR i IN 0 TO 12 GENERATE 
		wire_w_lg_doRR_pipe124w(i) <= doRR_pipe AND squarerIn1(i);
	END GENERATE loop149;
	loop150 : FOR i IN 0 TO 24 GENERATE 
		wire_w_lg_First_bit82w(i) <= First_bit AND man_above_half(i);
	END GENERATE loop150;
	loop151 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_small_flag214w(i) <= small_flag AND E_small(i);
	END GENERATE loop151;
	loop152 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_small_flag204w(i) <= small_flag AND wire_w203w(i);
	END GENERATE loop152;
	loop153 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_sR_pipe187w(i) <= sR_pipe1 AND wire_sub1_result(i);
	END GENERATE loop153;
	loop154 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_sR_pipe291w(i) <= sR_pipe2 AND wire_sub2_result(i);
	END GENERATE loop154;
	wire_w_lg_w_exp_data_range13w15w(0) <= wire_w_exp_data_range13w(0) AND wire_w_data_exp_is_ebiase_range6w(0);
	wire_w_lg_w_exp_data_range16w18w(0) <= wire_w_exp_data_range16w(0) AND wire_w_data_exp_is_ebiase_range14w(0);
	wire_w_lg_w_exp_data_range19w21w(0) <= wire_w_exp_data_range19w(0) AND wire_w_data_exp_is_ebiase_range17w(0);
	wire_w_lg_w_exp_data_range22w24w(0) <= wire_w_exp_data_range22w(0) AND wire_w_data_exp_is_ebiase_range20w(0);
	wire_w_lg_w_exp_data_range25w27w(0) <= wire_w_exp_data_range25w(0) AND wire_w_data_exp_is_ebiase_range23w(0);
	wire_w_lg_w_exp_data_range28w30w(0) <= wire_w_exp_data_range28w(0) AND wire_w_data_exp_is_ebiase_range26w(0);
	wire_w_lg_w_Log_g_range228w229w(0) <= wire_w_Log_g_range228w(0) AND wire_w_lg_w_Log_g_range226w227w(0);
	loop155 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_w_Log_small_range149w192w(i) <= wire_w_Log_small_range149w(0) AND wire_w_Log_small_range191w(i);
	END GENERATE loop155;
	loop156 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_w_Log_small_range150w197w(i) <= wire_w_Log_small_range150w(0) AND wire_w_Log_small_range196w(i);
	END GENERATE loop156;
	wire_w_lg_doRR111w(0) <= NOT doRR;
	wire_w_lg_doRR_pipe125w(0) <= NOT doRR_pipe;
	loop157 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_E_normal212w(i) <= NOT E_normal(i);
	END GENERATE loop157;
	wire_w_lg_exp_all_zero240w(0) <= NOT exp_all_zero;
	wire_w_lg_First_bit9w(0) <= NOT First_bit;
	wire_w_lg_input_is_one247w(0) <= NOT input_is_one;
	wire_w_lg_man_all_zero241w(0) <= NOT man_all_zero;
	wire_w_lg_small_flag206w(0) <= NOT small_flag;
	wire_w_lg_sR_pipe188w(0) <= NOT sR_pipe1;
	wire_w_lg_sR_pipe292w(0) <= NOT sR_pipe2;
	wire_w_lg_sR_pipe3179w(0) <= NOT sR_pipe3;
	wire_w_lg_w_E0_range38w39w(0) <= NOT wire_w_E0_range38w(0);
	wire_w_lg_w_E0_range42w43w(0) <= NOT wire_w_E0_range42w(0);
	wire_w_lg_w_E0_range46w47w(0) <= NOT wire_w_E0_range46w(0);
	wire_w_lg_w_E0_range50w51w(0) <= NOT wire_w_E0_range50w(0);
	wire_w_lg_w_E0_range54w55w(0) <= NOT wire_w_E0_range54w(0);
	wire_w_lg_w_E0_range58w59w(0) <= NOT wire_w_E0_range58w(0);
	wire_w_lg_w_E0_range62w63w(0) <= NOT wire_w_E0_range62w(0);
	wire_w_lg_w_E0_range66w67w(0) <= NOT wire_w_E0_range66w(0);
	wire_w_lg_w_exp_data_range31w33w(0) <= NOT wire_w_exp_data_range31w(0);
	wire_w_lg_w_Log_small_range149w154w(0) <= NOT wire_w_Log_small_range149w(0);
	wire_w_lg_w_Log_small_range150w198w(0) <= NOT wire_w_Log_small_range150w(0);
	wire_w_lg_w_lg_input_is_one247w248w(0) <= wire_w_lg_input_is_one247w(0) OR input_is_nan;
	wire_w_lg_w_lg_w_lg_input_is_zero244w245w246w(0) <= wire_w_lg_w_lg_input_is_zero244w245w(0) OR input_is_one;
	wire_w_lg_w_lg_input_is_zero244w245w(0) <= wire_w_lg_input_is_zero244w(0) OR input_is_nan;
	wire_w_lg_w_lg_sR254w255w(0) <= wire_w_lg_sR254w(0) OR input_is_nan;
	wire_w_lg_input_is_zero244w(0) <= input_is_zero OR input_is_infinity;
	wire_w_lg_sR254w(0) <= sR OR input_is_zero;
	wire_w_lg_w_Log_g_range220w221w(0) <= wire_w_Log_g_range220w(0) OR wire_w_sticky_range218w(0);
	wire_w_lg_w_Log_g_range223w224w(0) <= wire_w_Log_g_range223w(0) OR wire_w_sticky_range222w(0);
	wire_w_lg_w_Log_g_range226w227w(0) <= wire_w_Log_g_range226w(0) OR wire_w_sticky_range225w(0);
	wire_w_lg_w_Log_small_range150w155w(0) <= wire_w_Log_small_range150w(0) OR wire_w_lg_w_Log_small_range149w154w(0);
	wire_w_lg_w_Log_small_range150w151w(0) <= wire_w_Log_small_range150w(0) OR wire_w_Log_small_range149w(0);
	loop158 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_First_bit96w(i) <= First_bit XOR wire_w_Y0_range95w(i);
	END GENERATE loop158;
	absE <= (wire_w_lg_w_lg_sR_pipe292w93w OR wire_w_lg_sR_pipe291w);
	absELog2 <= absELog2_pipe_reg2;
	absELog2_pad <= ( absELog2 & "000000000000");
	absELog2_pipe <= wire_mult1_result;
	absZ0 <= absZ0_pipe_reg9;
	absZ0_pipe <= (wire_w_lg_w_lg_sR_pipe188w89w OR wire_w_lg_sR_pipe187w);
	absZ0s <= wire_Lshiftsmall_result(31 DOWNTO 20);
	absZ0s_pipe1 <= absZ0s_reg0;
	absZ0s_pipe2 <= absZ0s_pipe1_reg3;
	aclr <= '0';
	almostLog <= almostLog_pipe_reg2;
	almostLog_pipe <= wire_range_reduction_almostlog;
	clk_en <= '1';
	data_exp_is_ebiase <= ( wire_w_lg_w_lg_w_exp_data_range31w33w34w & wire_w_lg_w_exp_data_range28w30w & wire_w_lg_w_exp_data_range25w27w & wire_w_lg_w_exp_data_range22w24w & wire_w_lg_w_exp_data_range19w21w & wire_w_lg_w_exp_data_range16w18w & wire_w_lg_w_exp_data_range13w15w & exp_data(0));
	doRR <= Lshiftval(5);
	doRR_pipe <= doRR_reg1(0);
	E0 <= E0_pipe_reg9;
	E0_is_zero <= ( wire_w_lg_w_lg_w_E0_range66w67w68w & wire_w_lg_w_lg_w_E0_range62w63w64w & wire_w_lg_w_lg_w_E0_range58w59w60w & wire_w_lg_w_lg_w_E0_range54w55w56w & wire_w_lg_w_lg_w_E0_range50w51w52w & wire_w_lg_w_lg_w_E0_range46w47w48w & wire_w_lg_w_lg_w_E0_range42w43w44w & wire_w_lg_w_E0_range38w39w);
	E0_pipe <= wire_exp_biase_sub_result;
	E0_sub <= ( wire_w_lg_w_Log_small_range150w151w & wire_w_lg_w_Log_small_range150w155w);
	E0offset <= "10000110";
	E_normal <= E_normal_pipe_reg0;
	E_normal_pipe <= wire_lzc_norm_E_q(4 DOWNTO 0);
	E_small <= wire_sub5_result;
	EFR <= wire_add2_result;
	ER <= (wire_w_lg_w_lg_small_flag206w215w OR wire_w_lg_small_flag214w);
	exp_all_one <= wire_exp_nan_result;
	exp_all_zero <= wire_exp_zero_result;
	exp_biase <= ( "0111111" & wire_w_lg_First_bit9w);
	exp_data <= data(30 DOWNTO 23);
	exp_is_ebiase <= exp_is_ebiase_pipe_reg2(0);
	exp_is_ebiase_pipe <= data_exp_is_ebiase(7);
	First_bit <= man_data(22);
	input_is_infinity <= input_is_infinity_pipe_reg17(0);
	input_is_infinity_pipe <= (exp_all_one AND wire_w_lg_man_all_zero241w(0));
	input_is_nan <= input_is_nan_pipe_reg17(0);
	input_is_nan_pipe <= ((exp_all_one AND man_not_zero) OR sign_data_pipe);
	input_is_one <= input_is_one_pipe_reg17(0);
	input_is_one_pipe <= (exp_is_ebiase AND wire_w_lg_man_all_zero241w(0));
	input_is_zero <= input_is_zero_pipe_reg17(0);
	input_is_zero_pipe <= wire_w_lg_exp_all_zero240w(0);
	Log1p_normal <= wire_sub4_result;
	Log2 <= "101100010111001000011000000";
	Log_g <= (wire_w_lg_w_lg_small_flag206w207w OR wire_w_lg_small_flag204w);
	Log_normal <= wire_addsub2_result;
	Log_normal_normd <= Log_normal_normd_pipe_reg0;
	Log_normal_normd_pipe <= wire_lzc_norm_L_result(63 DOWNTO 17);
	Log_normal_pipe <= Log_normal_reg0;
	Log_small <= wire_addsub1_result;
	Log_small1 <= (wire_w_lg_w_lg_w_Log_small_range149w154w194w OR wire_w_lg_w_Log_small_range149w192w);
	Log_small2 <= (wire_w_lg_w_lg_w_Log_small_range150w198w199w OR wire_w_lg_w_Log_small_range150w197w);
	Log_small_normd <= Log_small_normd_pipe_reg1;
	Log_small_normd_pipe <= Log_small2;
	LogF_normal <= wire_add1_result;
	LogF_normal_pad <= ( LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal);
	Lshiftval <= wire_sub3_result;
	lzo <= lzo_pipe1_reg9;
	lzo_pipe1 <= (NOT wire_lzoc_q);
	lzo_pipe2 <= lzo_reg7;
	man_above_half <= ( "0" & "1" & man_data);
	man_all_zero <= wire_man_inf_result;
	man_below_half <= ( "1" & man_data & "0");
	man_data <= data(22 DOWNTO 0);
	man_not_zero <= wire_man_nan_result;
	nan <= input_is_nan;
	pfinal_s <= "01101";
	result <= ( wire_w_lg_w_lg_w_lg_sR254w255w256w & wire_mux_result0a_dataout);
	round <= wire_w_lg_w_Log_g_range228w229w(0);
	Rshiftval <= Lshiftval_reg3;
	sign_data <= data(31);
	sign_data_pipe <= sign_data_reg2(0);
	small_flag <= small_flag_pipe_reg9(0);
	small_flag_pipe <= (wire_w_lg_doRR111w(0) AND E0_is_zero(7));
	squarerIn <= (wire_w_lg_w_lg_doRR_pipe125w126w OR wire_w_lg_doRR_pipe124w);
	squarerIn0 <= ( absZ0s_pipe1 & "0");
	squarerIn1 <= Zfinal(25 DOWNTO 13);
	sR <= sR_pipe3_reg4(0);
	sR_pipe1 <= (NOT (data_exp_is_ebiase(7) OR exp_data(7)));
	sR_pipe2 <= sR_pipe1_reg9(0);
	sR_pipe3 <= sR_pipe2_reg5(0);
	sticky <= ( wire_w_lg_w_Log_g_range223w224w & wire_w_lg_w_Log_g_range220w221w & Log_g(0));
	wire_w203w <= ( Log_small_normd(25 DOWNTO 0) & "0");
	Y0 <= (wire_w_lg_w_lg_First_bit9w83w OR wire_w_lg_First_bit82w);
	Z2o2 <= Z2o2_pipe_reg0;
	Z2o2_pipe <= wire_squarer_result;
	Z2o2_small <= ( "0000000000000" & Z2o2_small_s & "00");
	Z2o2_small_s <= Z2o2_small_s_pipe_reg0;
	Z2o2_small_s_pipe <= wire_Rshiftsmall_result(31 DOWNTO 18);
	Z_small <= ( absZ0s_pipe2 & "00000000000000000");
	zero <= (input_is_one AND (NOT ((input_is_nan OR input_is_zero) OR input_is_infinity)));
	Zfinal <= wire_range_reduction_z;
	Zfinal_pipe <= Zfinal_reg1;
	wire_w_data_exp_is_ebiase_range6w(0) <= data_exp_is_ebiase(0);
	wire_w_data_exp_is_ebiase_range14w(0) <= data_exp_is_ebiase(1);
	wire_w_data_exp_is_ebiase_range17w(0) <= data_exp_is_ebiase(2);
	wire_w_data_exp_is_ebiase_range20w(0) <= data_exp_is_ebiase(3);
	wire_w_data_exp_is_ebiase_range23w(0) <= data_exp_is_ebiase(4);
	wire_w_data_exp_is_ebiase_range26w(0) <= data_exp_is_ebiase(5);
	wire_w_data_exp_is_ebiase_range29w(0) <= data_exp_is_ebiase(6);
	wire_w_E0_range38w(0) <= E0(0);
	wire_w_E0_range42w(0) <= E0(1);
	wire_w_E0_range46w(0) <= E0(2);
	wire_w_E0_range50w(0) <= E0(3);
	wire_w_E0_range54w(0) <= E0(4);
	wire_w_E0_range58w(0) <= E0(5);
	wire_w_E0_range62w(0) <= E0(6);
	wire_w_E0_range66w(0) <= E0(7);
	wire_w_E0_is_zero_range40w(0) <= E0_is_zero(0);
	wire_w_E0_is_zero_range45w(0) <= E0_is_zero(1);
	wire_w_E0_is_zero_range49w(0) <= E0_is_zero(2);
	wire_w_E0_is_zero_range53w(0) <= E0_is_zero(3);
	wire_w_E0_is_zero_range57w(0) <= E0_is_zero(4);
	wire_w_E0_is_zero_range61w(0) <= E0_is_zero(5);
	wire_w_E0_is_zero_range65w(0) <= E0_is_zero(6);
	wire_w_exp_data_range13w(0) <= exp_data(1);
	wire_w_exp_data_range16w(0) <= exp_data(2);
	wire_w_exp_data_range19w(0) <= exp_data(3);
	wire_w_exp_data_range22w(0) <= exp_data(4);
	wire_w_exp_data_range25w(0) <= exp_data(5);
	wire_w_exp_data_range28w(0) <= exp_data(6);
	wire_w_exp_data_range31w(0) <= exp_data(7);
	wire_w_Log_g_range220w(0) <= Log_g(1);
	wire_w_Log_g_range223w(0) <= Log_g(2);
	wire_w_Log_g_range228w(0) <= Log_g(3);
	wire_w_Log_g_range226w(0) <= Log_g(4);
	wire_w_Log_normal_normd_range205w <= Log_normal_normd(45 DOWNTO 19);
	wire_w_Log_small_range193w <= Log_small(26 DOWNTO 0);
	wire_w_Log_small_range191w <= Log_small(27 DOWNTO 1);
	wire_w_Log_small_range149w(0) <= Log_small(27);
	wire_w_Log_small_range196w <= Log_small(28 DOWNTO 2);
	wire_w_Log_small_range150w(0) <= Log_small(28);
	wire_w_sticky_range218w(0) <= sticky(0);
	wire_w_sticky_range222w(0) <= sticky(1);
	wire_w_sticky_range225w(0) <= sticky(2);
	wire_w_Y0_range86w <= Y0(11 DOWNTO 0);
	wire_w_Y0_range95w <= Y0(23 DOWNTO 1);
	wire_Lshiftsmall_data <= ( absZ0 & "00000000000000000000");
	Lshiftsmall :  fplog_altbarrel_shift_itd
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_Lshiftsmall_data,
		distance => Lshiftval(4 DOWNTO 0),
		result => wire_Lshiftsmall_result
	  );
	wire_lzc_norm_L_data <= ( Log_normal_pipe & "00000000000000000");
	wire_lzc_norm_L_distance <= wire_lzc_norm_E_w_lg_q189w;
	loop159 : FOR i IN 0 TO 5 GENERATE 
		wire_lzc_norm_E_w_lg_q189w(i) <= NOT wire_lzc_norm_E_q(i);
	END GENERATE loop159;
	lzc_norm_L :  fplog_altbarrel_shift_qab
	  PORT MAP ( 
		data => wire_lzc_norm_L_data,
		distance => wire_lzc_norm_L_distance,
		result => wire_lzc_norm_L_result
	  );
	wire_Rshiftsmall_data <= ( Z2o2 & "000000000000000000");
	Rshiftsmall :  fplog_altbarrel_shift_51e
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_Rshiftsmall_data,
		distance => Rshiftval(4 DOWNTO 0),
		result => wire_Rshiftsmall_result
	  );
	exp_nan :  fplog_altfp_log_and_or_h9b
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => exp_data,
		result => wire_exp_nan_result
	  );
	exp_zero :  fplog_altfp_log_and_or_v6b
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => exp_data,
		result => wire_exp_zero_result
	  );
	man_inf :  fplog_altfp_log_and_or_c8b
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => man_data,
		result => wire_man_inf_result
	  );
	man_nan :  fplog_altfp_log_and_or_c8b
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => man_data,
		result => wire_man_nan_result
	  );
	wire_add1_dataa <= ( "0000000000000" & Log1p_normal);
	add1 :  fplog_altfp_log_csa_s0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_add1_dataa,
		datab => almostLog,
		result => wire_add1_result
	  );
	wire_add2_dataa <= ( ER & Log_g(26 DOWNTO 4));
	wire_add2_datab <= ( "000000000000000000000000000000" & round);
	add2 :  fplog_altfp_log_csa_k0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_add2_dataa,
		datab => wire_add2_datab,
		result => wire_add2_result
	  );
	exp_biase_sub :  fplog_altfp_log_csa_0nc
	  PORT MAP ( 
		dataa => exp_data,
		datab => exp_biase,
		result => wire_exp_biase_sub_result
	  );
	wire_sub1_dataa <= (OTHERS => '0');
	sub1 :  fplog_altfp_log_csa_d4b
	  PORT MAP ( 
		dataa => wire_sub1_dataa,
		datab => Y0(11 DOWNTO 0),
		result => wire_sub1_result
	  );
	wire_sub2_dataa <= (OTHERS => '0');
	sub2 :  fplog_altfp_log_csa_0nc
	  PORT MAP ( 
		dataa => wire_sub2_dataa,
		datab => E0,
		result => wire_sub2_result
	  );
	wire_sub3_dataa <= ( "0" & lzo);
	wire_sub3_datab <= ( "0" & pfinal_s);
	sub3 :  fplog_altfp_log_csa_umc
	  PORT MAP ( 
		dataa => wire_sub3_dataa,
		datab => wire_sub3_datab,
		result => wire_sub3_result
	  );
	wire_sub4_datab <= ( "00000000000000" & Z2o2(13 DOWNTO 2));
	sub4 :  fplog_altfp_log_csa_nlf
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => Zfinal_pipe,
		datab => wire_sub4_datab,
		result => wire_sub4_result
	  );
	wire_sub5_dataa <= ( "0" & "11111" & E0_sub);
	wire_sub5_datab <= ( "000" & lzo_pipe2);
	sub5 :  fplog_altfp_log_csa_8kf
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_sub5_dataa,
		datab => wire_sub5_datab,
		result => wire_sub5_result
	  );
	wire_sub6_datab <= ( "000" & wire_w_lg_E_normal212w);
	sub6 :  fplog_altfp_log_csa_0nc
	  PORT MAP ( 
		dataa => E0offset,
		datab => wire_sub6_datab,
		result => wire_sub6_result
	  );
	range_reduction :  fplog_range_reduction_uqd
	  PORT MAP ( 
		a0_in => man_data(22 DOWNTO 18),
		aclr => aclr,
		almostlog => wire_range_reduction_almostlog,
		clk_en => clk_en,
		clock => clock,
		y0_in => Y0,
		z => wire_range_reduction_z
	  );
	wire_lzc_norm_E_data <= ( Log_normal & "00000000000000001");
	lzc_norm_E :  fplog_altpriority_encoder_uja
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_lzc_norm_E_data,
		q => wire_lzc_norm_E_q
	  );
	wire_lzoc_data <= ( wire_w_lg_First_bit96w & "000000001");
	lzoc :  fplog_altpriority_encoder_q08
	  PORT MAP ( 
		data => wire_lzoc_data,
		q => wire_lzoc_q
	  );
	squarer :  altsquare
	  GENERIC MAP (
		DATA_WIDTH => 13,
		PIPELINE => 1,
		REPRESENTATION => "UNSIGNED",
		RESULT_ALIGNMENT => "MSB",
		RESULT_WIDTH => 14
	  )
	  PORT MAP ( 
		aclr => aclr,
		clock => clock,
		data => squarerIn,
		ena => clk_en,
		result => wire_squarer_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absELog2_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absELog2_pipe_reg0 <= absELog2_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absELog2_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absELog2_pipe_reg1 <= absELog2_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absELog2_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absELog2_pipe_reg2 <= absELog2_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg0 <= absZ0_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg1 <= absZ0_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg2 <= absZ0_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg3 <= absZ0_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg4 <= absZ0_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg5 <= absZ0_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg6 <= absZ0_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg7 <= absZ0_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg8 <= absZ0_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg9 <= absZ0_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0s_pipe1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0s_pipe1_reg0 <= absZ0s_pipe1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0s_pipe1_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0s_pipe1_reg1 <= absZ0s_pipe1_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0s_pipe1_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0s_pipe1_reg2 <= absZ0s_pipe1_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0s_pipe1_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0s_pipe1_reg3 <= absZ0s_pipe1_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0s_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0s_reg0 <= absZ0s;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN almostLog_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN almostLog_pipe_reg0 <= almostLog_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN almostLog_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN almostLog_pipe_reg1 <= almostLog_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN almostLog_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN almostLog_pipe_reg2 <= almostLog_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN doRR_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN doRR_reg0(0) <= doRR;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN doRR_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN doRR_reg1 <= doRR_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg0 <= E0_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg1 <= E0_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg2 <= E0_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg3 <= E0_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg4 <= E0_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg5 <= E0_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg6 <= E0_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg7 <= E0_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg8 <= E0_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg9 <= E0_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E_normal_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E_normal_pipe_reg0 <= E_normal_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_is_ebiase_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_is_ebiase_pipe_reg0(0) <= exp_is_ebiase_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_is_ebiase_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_is_ebiase_pipe_reg1 <= exp_is_ebiase_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_is_ebiase_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_is_ebiase_pipe_reg2 <= exp_is_ebiase_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg0(0) <= input_is_infinity_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg1 <= input_is_infinity_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg10 <= input_is_infinity_pipe_reg9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg11 <= input_is_infinity_pipe_reg10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg12 <= input_is_infinity_pipe_reg11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg13 <= input_is_infinity_pipe_reg12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg14 <= input_is_infinity_pipe_reg13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg15 <= input_is_infinity_pipe_reg14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg16 <= input_is_infinity_pipe_reg15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg17 <= input_is_infinity_pipe_reg16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg2 <= input_is_infinity_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg3 <= input_is_infinity_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg4 <= input_is_infinity_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg5 <= input_is_infinity_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg6 <= input_is_infinity_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg7 <= input_is_infinity_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg8 <= input_is_infinity_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg9 <= input_is_infinity_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg0(0) <= input_is_nan_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg1 <= input_is_nan_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg10 <= input_is_nan_pipe_reg9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg11 <= input_is_nan_pipe_reg10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg12 <= input_is_nan_pipe_reg11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg13 <= input_is_nan_pipe_reg12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg14 <= input_is_nan_pipe_reg13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg15 <= input_is_nan_pipe_reg14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg16 <= input_is_nan_pipe_reg15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg17 <= input_is_nan_pipe_reg16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg2 <= input_is_nan_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg3 <= input_is_nan_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg4 <= input_is_nan_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg5 <= input_is_nan_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg6 <= input_is_nan_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg7 <= input_is_nan_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg8 <= input_is_nan_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg9 <= input_is_nan_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg0(0) <= input_is_one_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg1 <= input_is_one_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg10 <= input_is_one_pipe_reg9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg11 <= input_is_one_pipe_reg10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg12 <= input_is_one_pipe_reg11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg13 <= input_is_one_pipe_reg12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg14 <= input_is_one_pipe_reg13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg15 <= input_is_one_pipe_reg14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg16 <= input_is_one_pipe_reg15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg17 <= input_is_one_pipe_reg16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg2 <= input_is_one_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg3 <= input_is_one_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg4 <= input_is_one_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg5 <= input_is_one_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg6 <= input_is_one_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg7 <= input_is_one_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg8 <= input_is_one_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg9 <= input_is_one_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg0(0) <= input_is_zero_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg1 <= input_is_zero_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg10 <= input_is_zero_pipe_reg9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg11 <= input_is_zero_pipe_reg10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg12 <= input_is_zero_pipe_reg11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg13 <= input_is_zero_pipe_reg12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg14 <= input_is_zero_pipe_reg13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg15 <= input_is_zero_pipe_reg14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg16 <= input_is_zero_pipe_reg15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg17 <= input_is_zero_pipe_reg16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg2 <= input_is_zero_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg3 <= input_is_zero_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg4 <= input_is_zero_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg5 <= input_is_zero_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg6 <= input_is_zero_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg7 <= input_is_zero_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg8 <= input_is_zero_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg9 <= input_is_zero_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Log_normal_normd_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Log_normal_normd_pipe_reg0 <= Log_normal_normd_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Log_normal_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Log_normal_reg0 <= Log_normal;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Log_small_normd_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Log_small_normd_pipe_reg0 <= Log_small_normd_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Log_small_normd_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Log_small_normd_pipe_reg1 <= Log_small_normd_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Lshiftval_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Lshiftval_reg0 <= Lshiftval;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Lshiftval_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Lshiftval_reg1 <= Lshiftval_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Lshiftval_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Lshiftval_reg2 <= Lshiftval_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Lshiftval_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Lshiftval_reg3 <= Lshiftval_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg0 <= lzo_pipe1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg1 <= lzo_pipe1_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg2 <= lzo_pipe1_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg3 <= lzo_pipe1_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg4 <= lzo_pipe1_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg5 <= lzo_pipe1_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg6 <= lzo_pipe1_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg7 <= lzo_pipe1_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg8 <= lzo_pipe1_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg9 <= lzo_pipe1_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg0 <= lzo;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg1 <= lzo_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg2 <= lzo_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg3 <= lzo_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg4 <= lzo_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg5 <= lzo_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg6 <= lzo_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg7 <= lzo_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_data_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_data_reg0(0) <= sign_data;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_data_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_data_reg1 <= sign_data_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_data_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_data_reg2 <= sign_data_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg0(0) <= small_flag_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg1 <= small_flag_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg2 <= small_flag_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg3 <= small_flag_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg4 <= small_flag_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg5 <= small_flag_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg6 <= small_flag_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg7 <= small_flag_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg8 <= small_flag_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg9 <= small_flag_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg0(0) <= sR_pipe1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg1 <= sR_pipe1_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg2 <= sR_pipe1_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg3 <= sR_pipe1_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg4 <= sR_pipe1_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg5 <= sR_pipe1_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg6 <= sR_pipe1_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg7 <= sR_pipe1_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg8 <= sR_pipe1_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg9 <= sR_pipe1_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg0(0) <= sR_pipe2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg1 <= sR_pipe2_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg2 <= sR_pipe2_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg3 <= sR_pipe2_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg4 <= sR_pipe2_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg5 <= sR_pipe2_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe3_reg0(0) <= sR_pipe3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe3_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe3_reg1 <= sR_pipe3_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe3_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe3_reg2 <= sR_pipe3_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe3_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe3_reg3 <= sR_pipe3_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe3_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe3_reg4 <= sR_pipe3_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Z2o2_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Z2o2_pipe_reg0 <= Z2o2_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Z2o2_small_s_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Z2o2_small_s_pipe_reg0 <= Z2o2_small_s_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Zfinal_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Zfinal_reg0 <= Zfinal;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Zfinal_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Zfinal_reg1 <= Zfinal_reg0;
			END IF;
		END IF;
	END PROCESS;
	addsub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 29
	  )
	  PORT MAP ( 
		add_sub => sR_pipe3,
		clock => clock,
		dataa => Z_small,
		datab => Z2o2_small,
		result => wire_addsub1_result
	  );
	wire_addsub2_add_sub <= wire_w_lg_sR_pipe3179w(0);
	addsub2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 47
	  )
	  PORT MAP ( 
		add_sub => wire_addsub2_add_sub,
		clock => clock,
		dataa => absELog2_pad,
		datab => LogF_normal_pad,
		result => wire_addsub2_result
	  );
	mult1 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 8,
		LPM_WIDTHB => 27,
		LPM_WIDTHP => 35
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => absE,
		datab => Log2,
		result => wire_mult1_result
	  );
	wire_mux_result0a_dataout <= ( wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & input_is_nan & "0000000000000000000000") WHEN wire_w_lg_w_lg_w_lg_input_is_zero244w245w246w(0) = '1'  ELSE EFR;

 END RTL; --fplog_altfp_log_n6b
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY fplog IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		nan		: OUT STD_LOGIC ;
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		zero		: OUT STD_LOGIC 
	);
END fplog;


ARCHITECTURE RTL OF fplog IS

	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC ;



	COMPONENT fplog_altfp_log_n6b
	PORT (
			clock	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			nan	: OUT STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			zero	: OUT STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	nan    <= sub_wire0;
	result    <= sub_wire1(31 DOWNTO 0);
	zero    <= sub_wire2;

	fplog_altfp_log_n6b_component : fplog_altfp_log_n6b
	PORT MAP (
		clock => clock,
		data => data,
		nan => sub_wire0,
		result => sub_wire1,
		zero => sub_wire2
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_log"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "21"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: data 0 0 32 0 INPUT NODEFVAL "data[31..0]"
-- Retrieval info: CONNECT: @data 0 0 32 0 data 0 0 32 0
-- Retrieval info: USED_PORT: nan 0 0 0 0 OUTPUT NODEFVAL "nan"
-- Retrieval info: CONNECT: nan 0 0 0 0 @nan 0 0 0 0
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: USED_PORT: zero 0 0 0 0 OUTPUT NODEFVAL "zero"
-- Retrieval info: CONNECT: zero 0 0 0 0 @zero 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL fplog.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fplog.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fplog.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fplog_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fplog.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fplog.cmp TRUE TRUE
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX NUMERIC "1"
-- Retrieval info: LIB_FILE: lpm
