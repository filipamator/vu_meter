library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


entity fake_dac is
port (
        clock       : in STD_LOGIC;
        reset       : in STD_LOGIC;
        data_out    : out STD_LOGIC_VECTOR(15 downto 0);
        data_out_en : out STD_LOGIC
);
end fake_dac;


architecture Behavioral of fake_dac is


component gen48khz is
generic (
		CLKCOUNTER	: natural := 1000
);
port (
		clock 	: in std_logic;
		reset_n	: in std_logic;
		enable	: out std_logic
);
end component gen48khz;


signal counter      : integer;
signal sample_addr : integer range 0 to 8191;
signal sample_value  : STD_LOGIC_VECTOR(15 downto 0);

signal tick,reset_n : STD_LOGIC;

begin

reset_n <= not reset;

gen48khz_i1 : gen48khz
generic map (
		CLKCOUNTER  => 1000 -- 1000
)
port map (
		clock       => clock,
		reset_n     => reset_n,
		enable      => tick
);


process (clock,reset) 
begin
    if reset='1' then
        sample_addr <= 0;
    elsif clock='1' and clock'event then
        if tick='1' then
            data_out <= sample_value;
            data_out_en <= '1';
            if sample_addr=8191 then
                sample_addr <= 0;
            else
                sample_addr <= sample_addr + 1;
            end if;
        else
            data_out_en <= '0';
        end if;
    end if;
end process;


with sample_addr select sample_value <=
"0000000000000000" when 0,
"0011001011000110" when 1,
"0011110111010001" when 2,
"0001100001111101" when 3,
"1110000000000001" when 4,
"1100000010001101" when 5,
"1101001010111111" when 6,
"0000100001011010" when 7,
"0011011101101100" when 8,
"0011101100100000" when 9,
"0001000010010000" when 10,
"1101100100001011" when 11,
"1100000000000001" when 12,
"1101100100001011" when 13,
"0001000010010000" when 14,
"0011101100100000" when 15,
"0011011101101100" when 16,
"0000100001011010" when 17,
"1101001010111111" when 18,
"1100000010001101" when 19,
"1110000000000000" when 20,
"0001100001111101" when 21,
"0011110111010001" when 22,
"0011001011000110" when 23,
"0000000000000000" when 24,
"1100110100111010" when 25,
"1100001000101111" when 26,
"1110011110000011" when 27,
"0001111111111111" when 28,
"0011111101110011" when 29,
"0010110101000001" when 30,
"1111011110100110" when 31,
"1100100010010100" when 32,
"1100010011100000" when 33,
"1110111101110000" when 34,
"0010011011110101" when 35,
"0011111111111111" when 36,
"0010011011110110" when 37,
"1110111101110000" when 38,
"1100010011100000" when 39,
"1100100010010011" when 40,
"1111011110100110" when 41,
"0010110101000001" when 42,
"0011111101110011" when 43,
"0010000000000000" when 44,
"1110011110000011" when 45,
"1100001000101111" when 46,
"1100110100111010" when 47,
"0000000000000000" when 48,
"0011001011000110" when 49,
"0011110111010001" when 50,
"0001100001111110" when 51,
"1110000000000001" when 52,
"1100000010001101" when 53,
"1101001010111111" when 54,
"0000100001011010" when 55,
"0011011101101100" when 56,
"0011101100100000" when 57,
"0001000010010000" when 58,
"1101100100001011" when 59,
"1100000000000001" when 60,
"1101100100001010" when 61,
"0001000010010000" when 62,
"0011101100100000" when 63,
"0011011101101101" when 64,
"0000100001011010" when 65,
"1101001010111111" when 66,
"1100000010001101" when 67,
"1110000000000000" when 68,
"0001100001111101" when 69,
"0011110111010001" when 70,
"0011001011000110" when 71,
"0000000000000000" when 72,
"1100110100111010" when 73,
"1100001000101111" when 74,
"1110011110000010" when 75,
"0001111111111111" when 76,
"0011111101110011" when 77,
"0010110101000001" when 78,
"1111011110100110" when 79,
"1100100010010100" when 80,
"1100010011100000" when 81,
"1110111101110000" when 82,
"0010011011110101" when 83,
"0011111111111111" when 84,
"0010011011110110" when 85,
"1110111101110000" when 86,
"1100010011100000" when 87,
"1100100010010011" when 88,
"1111011110100110" when 89,
"0010110101000001" when 90,
"0011111101110011" when 91,
"0010000000000000" when 92,
"1110011110000011" when 93,
"1100001000101111" when 94,
"1100110100111010" when 95,
"0000000000000000" when 96,
"0011001011000110" when 97,
"0011110111010001" when 98,
"0001100001111110" when 99,
"1110000000000001" when 100,
"1100000010001101" when 101,
"1101001010111111" when 102,
"0000100001011010" when 103,
"0011011101101100" when 104,
"0011101100100000" when 105,
"0001000010010000" when 106,
"1101100100001011" when 107,
"1100000000000001" when 108,
"1101100100001010" when 109,
"0001000010010000" when 110,
"0011101100100000" when 111,
"0011011101101101" when 112,
"0000100001011010" when 113,
"1101001011000000" when 114,
"1100000010001101" when 115,
"1110000000000000" when 116,
"0001100001111101" when 117,
"0011110111010001" when 118,
"0011001011000110" when 119,
"0000000000000000" when 120,
"1100110100111010" when 121,
"1100001000101111" when 122,
"1110011110000010" when 123,
"0001111111111111" when 124,
"0011111101110011" when 125,
"0010110101000001" when 126,
"1111011110100110" when 127,
"1100100010010100" when 128,
"1100010011100000" when 129,
"1110111101110000" when 130,
"0010011011110101" when 131,
"0011111111111111" when 132,
"0010011011110110" when 133,
"1110111101110000" when 134,
"1100010011100000" when 135,
"1100100010010011" when 136,
"1111011110100110" when 137,
"0010110101000000" when 138,
"0011111101110011" when 139,
"0010000000000000" when 140,
"1110011110000011" when 141,
"1100001000101111" when 142,
"1100110100111010" when 143,
"0000000000000000" when 144,
"0011001011000110" when 145,
"0011110111010001" when 146,
"0001100001111110" when 147,
"1110000000000001" when 148,
"1100000010001101" when 149,
"1101001010111111" when 150,
"0000100001011010" when 151,
"0011011101101100" when 152,
"0011101100100001" when 153,
"0001000010010000" when 154,
"1101100100001011" when 155,
"1100000000000001" when 156,
"1101100100001010" when 157,
"0001000010010000" when 158,
"0011101100100000" when 159,
"0011011101101101" when 160,
"0000100001011011" when 161,
"1101001011000000" when 162,
"1100000010001101" when 163,
"1110000000000000" when 164,
"0001100001111101" when 165,
"0011110111010001" when 166,
"0011001011000110" when 167,
"0000000000000000" when 168,
"1100110100111011" when 169,
"1100001000101111" when 170,
"1110011110000010" when 171,
"0001111111111111" when 172,
"0011111101110011" when 173,
"0010110101000001" when 174,
"1111011110100111" when 175,
"1100100010010100" when 176,
"1100010011011111" when 177,
"1110111101101111" when 178,
"0010011011110101" when 179,
"0011111111111111" when 180,
"0010011011110110" when 181,
"1110111101110001" when 182,
"1100010011100000" when 183,
"1100100010010011" when 184,
"1111011110100101" when 185,
"0010110101000000" when 186,
"0011111101110011" when 187,
"0010000000000000" when 188,
"1110011110000011" when 189,
"1100001000101111" when 190,
"1100110100111010" when 191,
"0000000000000000" when 192,
"0011001011000101" when 193,
"0011110111010001" when 194,
"0001100001111110" when 195,
"1110000000000001" when 196,
"1100000010001101" when 197,
"1101001010111111" when 198,
"0000100001011001" when 199,
"0011011101101100" when 200,
"0011101100100001" when 201,
"0001000010010001" when 202,
"1101100100001011" when 203,
"1100000000000001" when 204,
"1101100100001010" when 205,
"0001000010001111" when 206,
"0011101100100000" when 207,
"0011011101101101" when 208,
"0000100001011011" when 209,
"1101001011000000" when 210,
"1100000010001101" when 211,
"1110000000000000" when 212,
"0001100001111101" when 213,
"0011110111010001" when 214,
"0011001011000110" when 215,
"0000000000000000" when 216,
"1100110100111011" when 217,
"1100001000101111" when 218,
"1110011110000010" when 219,
"0001111111111111" when 220,
"0011111101110011" when 221,
"0010110101000001" when 222,
"1111011110100111" when 223,
"1100100010010100" when 224,
"1100010011011111" when 225,
"1110111101101111" when 226,
"0010011011110101" when 227,
"0011111111111111" when 228,
"0010011011110110" when 229,
"1110111101110001" when 230,
"1100010011100000" when 231,
"1100100010010011" when 232,
"1111011110100101" when 233,
"0010110101000000" when 234,
"0011111101110011" when 235,
"0010000000000000" when 236,
"1110011110000011" when 237,
"1100001000101111" when 238,
"1100110100111010" when 239,
"0000000000000000" when 240,
"0011001011000101" when 241,
"0011110111010001" when 242,
"0001100001111110" when 243,
"1110000000000001" when 244,
"1100000010001101" when 245,
"1101001010111111" when 246,
"0000100001011001" when 247,
"0011011101101100" when 248,
"0011101100100001" when 249,
"0001000010010001" when 250,
"1101100100001011" when 251,
"1100000000000001" when 252,
"1101100100001010" when 253,
"0001000010001111" when 254,
"0011101100100000" when 255,
"0011011101101101" when 256,
"0000100001011011" when 257,
"1101001011000000" when 258,
"1100000010001101" when 259,
"1110000000000000" when 260,
"0001100001111101" when 261,
"0011110111010001" when 262,
"0011001011000110" when 263,
"0000000000000000" when 264,
"1100110100111011" when 265,
"1100001000101111" when 266,
"1110011110000010" when 267,
"0001111111111111" when 268,
"0011111101110011" when 269,
"0010110101000001" when 270,
"1111011110100111" when 271,
"1100100010010100" when 272,
"1100010011011111" when 273,
"1110111101101111" when 274,
"0010011011110101" when 275,
"0011111111111111" when 276,
"0010011011110110" when 277,
"1110111101110001" when 278,
"1100010011100000" when 279,
"1100100010010011" when 280,
"1111011110100101" when 281,
"0010110101000000" when 282,
"0011111101110011" when 283,
"0010000000000000" when 284,
"1110011110000011" when 285,
"1100001000101111" when 286,
"1100110100111010" when 287,
"0000000000000000" when 288,
"0011001011000101" when 289,
"0011110111010001" when 290,
"0001100001111110" when 291,
"1110000000000001" when 292,
"1100000010001101" when 293,
"1101001010111111" when 294,
"0000100001011001" when 295,
"0011011101101100" when 296,
"0011101100100001" when 297,
"0001000010010001" when 298,
"1101100100001011" when 299,
"1100000000000001" when 300,
"1101100100001010" when 301,
"0001000010001111" when 302,
"0011101100100000" when 303,
"0011011101101101" when 304,
"0000100001011011" when 305,
"1101001011000000" when 306,
"1100000010001101" when 307,
"1110000000000000" when 308,
"0001100001111100" when 309,
"0011110111010001" when 310,
"0011001011000110" when 311,
"0000000000000000" when 312,
"1100110100111011" when 313,
"1100001000101111" when 314,
"1110011110000010" when 315,
"0001111111111111" when 316,
"0011111101110011" when 317,
"0010110101000001" when 318,
"1111011110100111" when 319,
"1100100010010100" when 320,
"1100010011011111" when 321,
"1110111101101111" when 322,
"0010011011110101" when 323,
"0011111111111111" when 324,
"0010011011110110" when 325,
"1110111101110001" when 326,
"1100010011100000" when 327,
"1100100010010011" when 328,
"1111011110100101" when 329,
"0010110101000000" when 330,
"0011111101110011" when 331,
"0010000000000000" when 332,
"1110011110000100" when 333,
"1100001000101111" when 334,
"1100110100111010" when 335,
"1111111111111111" when 336,
"0011001011000101" when 337,
"0011110111010010" when 338,
"0001100001111110" when 339,
"1110000000000001" when 340,
"1100000010001101" when 341,
"1101001010111111" when 342,
"0000100001011001" when 343,
"0011011101101100" when 344,
"0011101100100001" when 345,
"0001000010010001" when 346,
"1101100100001011" when 347,
"1100000000000001" when 348,
"1101100100001010" when 349,
"0001000010001111" when 350,
"0011101100100000" when 351,
"0011011101101101" when 352,
"0000100001011011" when 353,
"1101001011000000" when 354,
"1100000010001101" when 355,
"1110000000000000" when 356,
"0001100001111100" when 357,
"0011110111010001" when 358,
"0011001011000110" when 359,
"0000000000000001" when 360,
"1100110100111011" when 361,
"1100001000101110" when 362,
"1110011110000010" when 363,
"0001111111111111" when 364,
"0011111101110011" when 365,
"0010110101000010" when 366,
"1111011110100111" when 367,
"1100100010010100" when 368,
"1100010011011111" when 369,
"1110111101101111" when 370,
"0010011011110101" when 371,
"0011111111111111" when 372,
"0010011011110110" when 373,
"1110111101110001" when 374,
"1100010011100000" when 375,
"1100100010010011" when 376,
"1111011110100101" when 377,
"0010110101000000" when 378,
"0011111101110011" when 379,
"0010000000000001" when 380,
"1110011110000100" when 381,
"1100001000101111" when 382,
"1100110100111001" when 383,
"1111111111111111" when 384,
"0011001011000101" when 385,
"0011110111010010" when 386,
"0001100001111111" when 387,
"1110000000000010" when 388,
"1100000010001101" when 389,
"1101001010111110" when 390,
"0000100001011001" when 391,
"0011011101101100" when 392,
"0011101100100001" when 393,
"0001000010010001" when 394,
"1101100100001100" when 395,
"1100000000000001" when 396,
"1101100100001010" when 397,
"0001000010001111" when 398,
"0011101100100000" when 399,
"0011011101101101" when 400,
"0000100001011011" when 401,
"1101001011000000" when 402,
"1100000010001101" when 403,
"1101111111111111" when 404,
"0001100001111100" when 405,
"0011110111010001" when 406,
"0011001011000111" when 407,
"0000000000000001" when 408,
"1100110100111011" when 409,
"1100001000101110" when 410,
"1110011110000001" when 411,
"0001111111111110" when 412,
"0011111101110011" when 413,
"0010110101000010" when 414,
"1111011110100111" when 415,
"1100100010010100" when 416,
"1100010011011111" when 417,
"1110111101101111" when 418,
"0010011011110100" when 419,
"0011111111111111" when 420,
"0010011011110110" when 421,
"1110111101110001" when 422,
"1100010011100000" when 423,
"1100100010010011" when 424,
"1111011110100101" when 425,
"0010110101000000" when 426,
"0011111101110100" when 427,
"0010000000000001" when 428,
"1110011110000100" when 429,
"1100001000101111" when 430,
"1100110100111001" when 431,
"1111111111111111" when 432,
"0011001011000101" when 433,
"0011110111010010" when 434,
"0001100001111111" when 435,
"1110000000000010" when 436,
"1100000010001101" when 437,
"1101001010111110" when 438,
"0000100001011001" when 439,
"0011011101101100" when 440,
"0011101100100001" when 441,
"0001000010010001" when 442,
"1101100100001100" when 443,
"1100000000000001" when 444,
"1101100100001001" when 445,
"0001000010001111" when 446,
"0011101100100000" when 447,
"0011011101101101" when 448,
"0000100001011011" when 449,
"1101001011000000" when 450,
"1100000010001100" when 451,
"1101111111111111" when 452,
"0001100001111100" when 453,
"0011110111010001" when 454,
"0011001011000111" when 455,
"0000000000000001" when 456,
"1100110100111011" when 457,
"1100001000101110" when 458,
"1110011110000001" when 459,
"0001111111111110" when 460,
"0011111101110011" when 461,
"0010110101000010" when 462,
"1111011110100111" when 463,
"1100100010010100" when 464,
"1100010011011111" when 465,
"1110111101101111" when 466,
"0010011011110100" when 467,
"0011111111111111" when 468,
"0010011011110111" when 469,
"1110111101110001" when 470,
"1100010011100000" when 471,
"1100100010010011" when 472,
"1111011110100100" when 473,
"0010110101000000" when 474,
"0011111101110100" when 475,
"0010000000000001" when 476,
"1110011110000100" when 477,
"1100001000101111" when 478,
"1100110100111001" when 479,
"1111111111111111" when 480,
"0011001011000101" when 481,
"0011110111010010" when 482,
"0001100001111111" when 483,
"1110000000000010" when 484,
"1100000010001101" when 485,
"1101001010111110" when 486,
"0000100001011001" when 487,
"0011011101101100" when 488,
"0011101100100001" when 489,
"0001000010010001" when 490,
"1101100100001100" when 491,
"1100000000000001" when 492,
"1101100100001001" when 493,
"0001000010001111" when 494,
"0011101100100000" when 495,
"0011011101101101" when 496,
"0000100001011100" when 497,
"1101001011000000" when 498,
"1100000010001100" when 499,
"1101111111111111" when 500,
"0001100001111100" when 501,
"0011110111010001" when 502,
"0011001011000111" when 503,
"0000000000000001" when 504,
"1100110100111011" when 505,
"1100001000101110" when 506,
"1110011110000001" when 507,
"0001111111111110" when 508,
"0011111101110011" when 509,
"0010110101000010" when 510,
"1111011110101000" when 511,
"1100100010010100" when 512,
"1100010011011111" when 513,
"1110111101101110" when 514,
"0010011011110100" when 515,
"0011111111111111" when 516,
"0010011011110111" when 517,
"1110111101110010" when 518,
"1100010011100000" when 519,
"1100100010010011" when 520,
"1111011110100100" when 521,
"0010110101000000" when 522,
"0011111101110100" when 523,
"0010000000000001" when 524,
"1110011110000100" when 525,
"1100001000101111" when 526,
"1100110100111001" when 527,
"1111111111111111" when 528,
"0011001011000101" when 529,
"0011110111010010" when 530,
"0001100001111111" when 531,
"1110000000000010" when 532,
"1100000010001101" when 533,
"1101001010111110" when 534,
"0000100001011000" when 535,
"0011011101101100" when 536,
"0011101100100001" when 537,
"0001000010010010" when 538,
"1101100100001100" when 539,
"1100000000000001" when 540,
"1101100100001001" when 541,
"0001000010001110" when 542,
"0011101100100000" when 543,
"0011011101101101" when 544,
"0000100001011100" when 545,
"1101001011000000" when 546,
"1100000010001100" when 547,
"1101111111111111" when 548,
"0001100001111100" when 549,
"0011110111010001" when 550,
"0011001011000111" when 551,
"0000000000000001" when 552,
"1100110100111011" when 553,
"1100001000101110" when 554,
"1110011110000001" when 555,
"0001111111111110" when 556,
"0011111101110011" when 557,
"0010110101000010" when 558,
"1111011110101000" when 559,
"1100100010010100" when 560,
"1100010011011111" when 561,
"1110111101101110" when 562,
"0010011011110100" when 563,
"0011111111111111" when 564,
"0010011011110111" when 565,
"1110111101110010" when 566,
"1100010011100000" when 567,
"1100100010010011" when 568,
"1111011110100100" when 569,
"0010110100111111" when 570,
"0011111101110100" when 571,
"0010000000000001" when 572,
"1110011110000100" when 573,
"1100001000101111" when 574,
"1100110100111001" when 575,
"1111111111111111" when 576,
"0011001011000101" when 577,
"0011110111010010" when 578,
"0001100001111111" when 579,
"1110000000000010" when 580,
"1100000010001101" when 581,
"1101001010111110" when 582,
"0000100001011000" when 583,
"0011011101101100" when 584,
"0011101100100001" when 585,
"0001000010010010" when 586,
"1101100100001100" when 587,
"1100000000000001" when 588,
"1101100100001001" when 589,
"0001000010001110" when 590,
"0011101100100000" when 591,
"0011011101101101" when 592,
"0000100001011100" when 593,
"1101001011000001" when 594,
"1100000010001100" when 595,
"1101111111111111" when 596,
"0001100001111100" when 597,
"0011110111010001" when 598,
"0011001011000111" when 599,
"0000000000000001" when 600,
"1100110100111011" when 601,
"1100001000101110" when 602,
"1110011110000001" when 603,
"0001111111111110" when 604,
"0011111101110011" when 605,
"0010110101000010" when 606,
"1111011110101000" when 607,
"1100100010010100" when 608,
"1100010011011111" when 609,
"1110111101101110" when 610,
"0010011011110100" when 611,
"0011111111111111" when 612,
"0010011011110111" when 613,
"1110111101110010" when 614,
"1100010011100000" when 615,
"1100100010010011" when 616,
"1111011110100100" when 617,
"0010110100111111" when 618,
"0011111101110100" when 619,
"0010000000000001" when 620,
"1110011110000100" when 621,
"1100001000101111" when 622,
"1100110100111001" when 623,
"1111111111111111" when 624,
"0011001011000101" when 625,
"0011110111010010" when 626,
"0001100001111111" when 627,
"1110000000000010" when 628,
"1100000010001101" when 629,
"1101001010111110" when 630,
"0000100001011000" when 631,
"0011011101101011" when 632,
"0011101100100001" when 633,
"0001000010010010" when 634,
"1101100100001100" when 635,
"1100000000000001" when 636,
"1101100100001001" when 637,
"0001000010001110" when 638,
"0011101100100000" when 639,
"0011011101101101" when 640,
"0000100001011100" when 641,
"1101001011000001" when 642,
"1100000010001100" when 643,
"1101111111111111" when 644,
"0001100001111100" when 645,
"0011110111010001" when 646,
"0011001011000111" when 647,
"0000000000000010" when 648,
"1100110100111011" when 649,
"1100001000101110" when 650,
"1110011110000001" when 651,
"0001111111111110" when 652,
"0011111101110011" when 653,
"0010110101000010" when 654,
"1111011110101000" when 655,
"1100100010010101" when 656,
"1100010011011111" when 657,
"1110111101101110" when 658,
"0010011011110100" when 659,
"0011111111111111" when 660,
"0010011011110111" when 661,
"1110111101110010" when 662,
"1100010011100000" when 663,
"1100100010010011" when 664,
"1111011110100100" when 665,
"0010110100111111" when 666,
"0011111101110100" when 667,
"0010000000000001" when 668,
"1110011110000101" when 669,
"1100001000101111" when 670,
"1100110100111001" when 671,
"1111111111111110" when 672,
"0011001011000101" when 673,
"0011110111010010" when 674,
"0001100001111111" when 675,
"1110000000000010" when 676,
"1100000010001101" when 677,
"1101001010111110" when 678,
"0000100001011000" when 679,
"0011011101101011" when 680,
"0011101100100001" when 681,
"0001000010010010" when 682,
"1101100100001100" when 683,
"1100000000000001" when 684,
"1101100100001001" when 685,
"0001000010001110" when 686,
"0011101100100000" when 687,
"0011011101101110" when 688,
"0000100001011100" when 689,
"1101001011000001" when 690,
"1100000010001100" when 691,
"1101111111111111" when 692,
"0001100001111011" when 693,
"0011110111010001" when 694,
"0011001011000111" when 695,
"0000000000000010" when 696,
"1100110100111100" when 697,
"1100001000101110" when 698,
"1110011110000001" when 699,
"0001111111111110" when 700,
"0011111101110011" when 701,
"0010110101000010" when 702,
"1111011110101000" when 703,
"1100100010010101" when 704,
"1100010011011111" when 705,
"1110111101101110" when 706,
"0010011011110100" when 707,
"0011111111111111" when 708,
"0010011011110111" when 709,
"1110111101110010" when 710,
"1100010011100001" when 711,
"1100100010010010" when 712,
"1111011110100100" when 713,
"0010110100111111" when 714,
"0011111101110100" when 715,
"0010000000000001" when 716,
"1110011110000101" when 717,
"1100001000101111" when 718,
"1100110100111001" when 719,
"1111111111111110" when 720,
"0011001011000100" when 721,
"0011110111010010" when 722,
"0001100001111111" when 723,
"1110000000000010" when 724,
"1100000010001101" when 725,
"1101001010111110" when 726,
"0000100001011000" when 727,
"0011011101101011" when 728,
"0011101100100001" when 729,
"0001000010010010" when 730,
"1101100100001100" when 731,
"1100000000000001" when 732,
"1101100100001001" when 733,
"0001000010001110" when 734,
"0011101100011111" when 735,
"0011011101101110" when 736,
"0000100001011100" when 737,
"1101001011000001" when 738,
"1100000010001100" when 739,
"1101111111111110" when 740,
"0001100001111011" when 741,
"0011110111010001" when 742,
"0011001011000111" when 743,
"0000000000000010" when 744,
"1100110100111100" when 745,
"1100001000101110" when 746,
"1110011110000000" when 747,
"0001111111111101" when 748,
"0011111101110011" when 749,
"0010110101000010" when 750,
"1111011110101000" when 751,
"1100100010010101" when 752,
"1100010011011111" when 753,
"1110111101101110" when 754,
"0010011011110100" when 755,
"0011111111111111" when 756,
"0010011011110111" when 757,
"1110111101110010" when 758,
"1100010011100001" when 759,
"1100100010010010" when 760,
"1111011110100100" when 761,
"0010110100111111" when 762,
"0011111101110100" when 763,
"0010000000000010" when 764,
"1110011110000101" when 765,
"1100001000101111" when 766,
"1100110100111001" when 767,
"1111111111111110" when 768,
"0011001011000100" when 769,
"0011110111010010" when 770,
"0001100010000000" when 771,
"1110000000000011" when 772,
"1100000010001101" when 773,
"1101001010111110" when 774,
"0000100001011000" when 775,
"0011011101101011" when 776,
"0011101100100001" when 777,
"0001000010010010" when 778,
"1101100100001100" when 779,
"1100000000000001" when 780,
"1101100100001001" when 781,
"0001000010001110" when 782,
"0011101100011111" when 783,
"0011011101101110" when 784,
"0000100001011100" when 785,
"1101001011000001" when 786,
"1100000010001100" when 787,
"1101111111111110" when 788,
"0001100001111011" when 789,
"0011110111010001" when 790,
"0011001011000111" when 791,
"0000000000000010" when 792,
"1100110100111100" when 793,
"1100001000101110" when 794,
"1110011110000000" when 795,
"0001111111111101" when 796,
"0011111101110011" when 797,
"0010110101000010" when 798,
"1111011110101000" when 799,
"1100100010010101" when 800,
"1100010011011111" when 801,
"1110111101101110" when 802,
"0010011011110011" when 803,
"0011111111111111" when 804,
"0010011011110111" when 805,
"1110111101110010" when 806,
"1100010011100001" when 807,
"1100100010010010" when 808,
"1111011110100011" when 809,
"0010110100111111" when 810,
"0011111101110100" when 811,
"0010000000000010" when 812,
"1110011110000101" when 813,
"1100001000101111" when 814,
"1100110100111001" when 815,
"1111111111111110" when 816,
"0011001011000100" when 817,
"0011110111010010" when 818,
"0001100010000000" when 819,
"1110000000000011" when 820,
"1100000010001101" when 821,
"1101001010111101" when 822,
"0000100001010111" when 823,
"0011011101101011" when 824,
"0011101100100001" when 825,
"0001000010010010" when 826,
"1101100100001101" when 827,
"1100000000000001" when 828,
"1101100100001000" when 829,
"0001000010001101" when 830,
"0011101100011111" when 831,
"0011011101101110" when 832,
"0000100001011101" when 833,
"1101001011000001" when 834,
"1100000010001100" when 835,
"1101111111111110" when 836,
"0001100001111011" when 837,
"0011110111010001" when 838,
"0011001011000111" when 839,
"0000000000000010" when 840,
"1100110100111100" when 841,
"1100001000101110" when 842,
"1110011110000000" when 843,
"0001111111111101" when 844,
"0011111101110011" when 845,
"0010110101000011" when 846,
"1111011110101001" when 847,
"1100100010010101" when 848,
"1100010011011111" when 849,
"1110111101101101" when 850,
"0010011011110011" when 851,
"0011111111111111" when 852,
"0010011011111000" when 853,
"1110111101110011" when 854,
"1100010011100001" when 855,
"1100100010010010" when 856,
"1111011110100011" when 857,
"0010110100111111" when 858,
"0011111101110100" when 859,
"0010000000000010" when 860,
"1110011110000101" when 861,
"1100001000101111" when 862,
"1100110100111001" when 863,
"1111111111111110" when 864,
"0011001011000100" when 865,
"0011110111010010" when 866,
"0001100010000000" when 867,
"1110000000000011" when 868,
"1100000010001101" when 869,
"1101001010111101" when 870,
"0000100001010111" when 871,
"0011011101101011" when 872,
"0011101100100001" when 873,
"0001000010010011" when 874,
"1101100100001101" when 875,
"1100000000000001" when 876,
"1101100100001000" when 877,
"0001000010001101" when 878,
"0011101100011111" when 879,
"0011011101101110" when 880,
"0000100001011101" when 881,
"1101001011000001" when 882,
"1100000010001100" when 883,
"1101111111111110" when 884,
"0001100001111011" when 885,
"0011110111010001" when 886,
"0011001011000111" when 887,
"0000000000000010" when 888,
"1100110100111100" when 889,
"1100001000101110" when 890,
"1110011110000000" when 891,
"0001111111111101" when 892,
"0011111101110011" when 893,
"0010110101000011" when 894,
"1111011110101001" when 895,
"1100100010010101" when 896,
"1100010011011111" when 897,
"1110111101101101" when 898,
"0010011011110011" when 899,
"0011111111111111" when 900,
"0010011011111000" when 901,
"1110111101110011" when 902,
"1100010011100001" when 903,
"1100100010010010" when 904,
"1111011110100011" when 905,
"0010110100111111" when 906,
"0011111101110100" when 907,
"0010000000000010" when 908,
"1110011110000101" when 909,
"1100001000110000" when 910,
"1100110100111000" when 911,
"1111111111111110" when 912,
"0011001011000100" when 913,
"0011110111010010" when 914,
"0001100010000000" when 915,
"1110000000000011" when 916,
"1100000010001101" when 917,
"1101001010111101" when 918,
"0000100001010111" when 919,
"0011011101101011" when 920,
"0011101100100001" when 921,
"0001000010010011" when 922,
"1101100100001101" when 923,
"1100000000000001" when 924,
"1101100100001000" when 925,
"0001000010001101" when 926,
"0011101100011111" when 927,
"0011011101101110" when 928,
"0000100001011101" when 929,
"1101001011000001" when 930,
"1100000010001100" when 931,
"1101111111111110" when 932,
"0001100001111011" when 933,
"0011110111010000" when 934,
"0011001011001000" when 935,
"0000000000000010" when 936,
"1100110100111100" when 937,
"1100001000101110" when 938,
"1110011110000000" when 939,
"0001111111111101" when 940,
"0011111101110011" when 941,
"0010110101000011" when 942,
"1111011110101001" when 943,
"1100100010010101" when 944,
"1100010011011111" when 945,
"1110111101101101" when 946,
"0010011011110011" when 947,
"0011111111111111" when 948,
"0010011011111000" when 949,
"1110111101110011" when 950,
"1100010011100001" when 951,
"1100100010010010" when 952,
"1111011110100011" when 953,
"0010110100111111" when 954,
"0011111101110100" when 955,
"0010000000000010" when 956,
"1110011110000101" when 957,
"1100001000110000" when 958,
"1100110100111000" when 959,
"1111111111111110" when 960,
"0011001011000100" when 961,
"0011110111010010" when 962,
"0001100010000000" when 963,
"1110000000000011" when 964,
"1100000010001101" when 965,
"1101001010111101" when 966,
"0000100001010111" when 967,
"0011011101101011" when 968,
"0011101100100010" when 969,
"0001000010010011" when 970,
"1101100100001101" when 971,
"1100000000000001" when 972,
"1101100100001000" when 973,
"0001000010001101" when 974,
"0011101100011111" when 975,
"0011011101101110" when 976,
"0000100001011101" when 977,
"1101001011000001" when 978,
"1100000010001100" when 979,
"1101111111111110" when 980,
"0001100001111011" when 981,
"0011110111010000" when 982,
"0011001011001000" when 983,
"0000000000000011" when 984,
"1100110100111100" when 985,
"1100001000101110" when 986,
"1110011110000000" when 987,
"0001111111111101" when 988,
"0011111101110011" when 989,
"0010110101000011" when 990,
"1111011110101001" when 991,
"1100100010010101" when 992,
"1100010011011110" when 993,
"1110111101101101" when 994,
"0010011011110011" when 995,
"0011111111111111" when 996,
"0010011011111000" when 997,
"1110111101110011" when 998,
"1100010011100001" when 999,
"1100100010010010" when 1000,
"1111011110100011" when 1001,
"0010110100111111" when 1002,
"0011111101110100" when 1003,
"0010000000000010" when 1004,
"1110011110000110" when 1005,
"1100001000110000" when 1006,
"1100110100111000" when 1007,
"1111111111111101" when 1008,
"0011001011000100" when 1009,
"0011110111010010" when 1010,
"0001100010000000" when 1011,
"1110000000000011" when 1012,
"1100000010001101" when 1013,
"1101001010111101" when 1014,
"0000100001010111" when 1015,
"0011011101101011" when 1016,
"0011101100100010" when 1017,
"0001000010010011" when 1018,
"1101100100001101" when 1019,
"1100000000000001" when 1020,
"1101100100001000" when 1021,
"0001000010001101" when 1022,
"0011101100011111" when 1023,
"0011011101101110" when 1024,
"0000100001011101" when 1025,
"1101001011000010" when 1026,
"1100000010001100" when 1027,
"1101111111111110" when 1028,
"0001100001111010" when 1029,
"0011110111010000" when 1030,
"0011001011001000" when 1031,
"0000000000000011" when 1032,
"1100110100111100" when 1033,
"1100001000101110" when 1034,
"1110011110000000" when 1035,
"0001111111111101" when 1036,
"0011111101110011" when 1037,
"0010110101000011" when 1038,
"1111011110101001" when 1039,
"1100100010010101" when 1040,
"1100010011011110" when 1041,
"1110111101101101" when 1042,
"0010011011110011" when 1043,
"0011111111111111" when 1044,
"0010011011111000" when 1045,
"1110111101110011" when 1046,
"1100010011100001" when 1047,
"1100100010010010" when 1048,
"1111011110100011" when 1049,
"0010110100111110" when 1050,
"0011111101110100" when 1051,
"0010000000000010" when 1052,
"1110011110000110" when 1053,
"1100001000110000" when 1054,
"1100110100111000" when 1055,
"1111111111111101" when 1056,
"0011001011000100" when 1057,
"0011110111010010" when 1058,
"0001100010000000" when 1059,
"1110000000000011" when 1060,
"1100000010001101" when 1061,
"1101001010111101" when 1062,
"0000100001010111" when 1063,
"0011011101101011" when 1064,
"0011101100100010" when 1065,
"0001000010010011" when 1066,
"1101100100001101" when 1067,
"1100000000000001" when 1068,
"1101100100001000" when 1069,
"0001000010001101" when 1070,
"0011101100011111" when 1071,
"0011011101101110" when 1072,
"0000100001011101" when 1073,
"1101001011000010" when 1074,
"1100000010001100" when 1075,
"1101111111111110" when 1076,
"0001100001111010" when 1077,
"0011110111010000" when 1078,
"0011001011001000" when 1079,
"0000000000000011" when 1080,
"1100110100111100" when 1081,
"1100001000101110" when 1082,
"1110011101111111" when 1083,
"0001111111111101" when 1084,
"0011111101110011" when 1085,
"0010110101000011" when 1086,
"1111011110101001" when 1087,
"1100100010010101" when 1088,
"1100010011011110" when 1089,
"1110111101101101" when 1090,
"0010011011110011" when 1091,
"0011111111111111" when 1092,
"0010011011111000" when 1093,
"1110111101110011" when 1094,
"1100010011100001" when 1095,
"1100100010010010" when 1096,
"1111011110100011" when 1097,
"0010110100111110" when 1098,
"0011111101110100" when 1099,
"0010000000000010" when 1100,
"1110011110000110" when 1101,
"1100001000110000" when 1102,
"1100110100111000" when 1103,
"1111111111111101" when 1104,
"0011001011000100" when 1105,
"0011110111010010" when 1106,
"0001100010000001" when 1107,
"1110000000000011" when 1108,
"1100000010001101" when 1109,
"1101001010111101" when 1110,
"0000100001010111" when 1111,
"0011011101101011" when 1112,
"0011101100100010" when 1113,
"0001000010010011" when 1114,
"1101100100001101" when 1115,
"1100000000000001" when 1116,
"1101100100001000" when 1117,
"0001000010001101" when 1118,
"0011101100011111" when 1119,
"0011011101101110" when 1120,
"0000100001011110" when 1121,
"1101001011000010" when 1122,
"1100000010001100" when 1123,
"1101111111111101" when 1124,
"0001100001111010" when 1125,
"0011110111010000" when 1126,
"0011001011001000" when 1127,
"0000000000000011" when 1128,
"1100110100111100" when 1129,
"1100001000101110" when 1130,
"1110011101111111" when 1131,
"0001111111111100" when 1132,
"0011111101110011" when 1133,
"0010110101000011" when 1134,
"1111011110101001" when 1135,
"1100100010010101" when 1136,
"1100010011011110" when 1137,
"1110111101101101" when 1138,
"0010011011110011" when 1139,
"0011111111111111" when 1140,
"0010011011111000" when 1141,
"1110111101110011" when 1142,
"1100010011100001" when 1143,
"1100100010010010" when 1144,
"1111011110100010" when 1145,
"0010110100111110" when 1146,
"0011111101110100" when 1147,
"0010000000000011" when 1148,
"1110011110000110" when 1149,
"1100001000110000" when 1150,
"1100110100111000" when 1151,
"1111111111111101" when 1152,
"0011001011000100" when 1153,
"0011110111010010" when 1154,
"0001100010000001" when 1155,
"1110000000000100" when 1156,
"1100000010001101" when 1157,
"1101001010111101" when 1158,
"0000100001010110" when 1159,
"0011011101101011" when 1160,
"0011101100100010" when 1161,
"0001000010010011" when 1162,
"1101100100001101" when 1163,
"1100000000000001" when 1164,
"1101100100001000" when 1165,
"0001000010001100" when 1166,
"0011101100011111" when 1167,
"0011011101101110" when 1168,
"0000100001011110" when 1169,
"1101001011000010" when 1170,
"1100000010001100" when 1171,
"1101111111111101" when 1172,
"0001100001111010" when 1173,
"0011110111010000" when 1174,
"0011001011001000" when 1175,
"0000000000000011" when 1176,
"1100110100111100" when 1177,
"1100001000101110" when 1178,
"1110011101111111" when 1179,
"0001111111111100" when 1180,
"0011111101110011" when 1181,
"0010110101000011" when 1182,
"1111011110101010" when 1183,
"1100100010010101" when 1184,
"1100010011011110" when 1185,
"1110111101101100" when 1186,
"0010011011110011" when 1187,
"0011111111111111" when 1188,
"0010011011111000" when 1189,
"1110111101110100" when 1190,
"1100010011100001" when 1191,
"1100100010010010" when 1192,
"1111011110100010" when 1193,
"0010110100111110" when 1194,
"0011111101110100" when 1195,
"0010000000000011" when 1196,
"1110011110000110" when 1197,
"1100001000110000" when 1198,
"1100110100111000" when 1199,
"1111111111111101" when 1200,
"0011001011000100" when 1201,
"0011110111010010" when 1202,
"0001100010000001" when 1203,
"1110000000000100" when 1204,
"1100000010001101" when 1205,
"1101001010111101" when 1206,
"0000100001010110" when 1207,
"0011011101101011" when 1208,
"0011101100100010" when 1209,
"0001000010010100" when 1210,
"1101100100001110" when 1211,
"1100000000000001" when 1212,
"1101100100001000" when 1213,
"0001000010001100" when 1214,
"0011101100011111" when 1215,
"0011011101101110" when 1216,
"0000100001011110" when 1217,
"1101001011000010" when 1218,
"1100000010001100" when 1219,
"1101111111111101" when 1220,
"0001100001111010" when 1221,
"0011110111010000" when 1222,
"0011001011001000" when 1223,
"0000000000000011" when 1224,
"1100110100111101" when 1225,
"1100001000101110" when 1226,
"1110011101111111" when 1227,
"0001111111111100" when 1228,
"0011111101110011" when 1229,
"0010110101000011" when 1230,
"1111011110101010" when 1231,
"1100100010010101" when 1232,
"1100010011011110" when 1233,
"1110111101101100" when 1234,
"0010011011110010" when 1235,
"0011111111111111" when 1236,
"0010011011111001" when 1237,
"1110111101110100" when 1238,
"1100010011100001" when 1239,
"1100100010010010" when 1240,
"1111011110100010" when 1241,
"0010110100111110" when 1242,
"0011111101110100" when 1243,
"0010000000000011" when 1244,
"1110011110000110" when 1245,
"1100001000110000" when 1246,
"1100110100111000" when 1247,
"1111111111111101" when 1248,
"0011001011000011" when 1249,
"0011110111010010" when 1250,
"0001100010000001" when 1251,
"1110000000000100" when 1252,
"1100000010001101" when 1253,
"1101001010111100" when 1254,
"0000100001010110" when 1255,
"0011011101101010" when 1256,
"0011101100100010" when 1257,
"0001000010010100" when 1258,
"1101100100001110" when 1259,
"1100000000000001" when 1260,
"1101100100000111" when 1261,
"0001000010001100" when 1262,
"0011101100011111" when 1263,
"0011011101101110" when 1264,
"0000100001011110" when 1265,
"1101001011000010" when 1266,
"1100000010001100" when 1267,
"1101111111111101" when 1268,
"0001100001111010" when 1269,
"0011110111010000" when 1270,
"0011001011001000" when 1271,
"0000000000000011" when 1272,
"1100110100111101" when 1273,
"1100001000101110" when 1274,
"1110011101111111" when 1275,
"0001111111111100" when 1276,
"0011111101110011" when 1277,
"0010110101000100" when 1278,
"1111011110101010" when 1279,
"1100100010010110" when 1280,
"1100010011011110" when 1281,
"1110111101101100" when 1282,
"0010011011110010" when 1283,
"0011111111111111" when 1284,
"0010011011111001" when 1285,
"1110111101110100" when 1286,
"1100010011100001" when 1287,
"1100100010010010" when 1288,
"1111011110100010" when 1289,
"0010110100111110" when 1290,
"0011111101110100" when 1291,
"0010000000000011" when 1292,
"1110011110000110" when 1293,
"1100001000110000" when 1294,
"1100110100111000" when 1295,
"1111111111111100" when 1296,
"0011001011000011" when 1297,
"0011110111010010" when 1298,
"0001100010000001" when 1299,
"1110000000000100" when 1300,
"1100000010001101" when 1301,
"1101001010111100" when 1302,
"0000100001010110" when 1303,
"0011011101101010" when 1304,
"0011101100100010" when 1305,
"0001000010010100" when 1306,
"1101100100001110" when 1307,
"1100000000000001" when 1308,
"1101100100000111" when 1309,
"0001000010001100" when 1310,
"0011101100011111" when 1311,
"0011011101101111" when 1312,
"0000100001011110" when 1313,
"1101001011000010" when 1314,
"1100000010001100" when 1315,
"1101111111111101" when 1316,
"0001100001111010" when 1317,
"0011110111010000" when 1318,
"0011001011001000" when 1319,
"0000000000000100" when 1320,
"1100110100111101" when 1321,
"1100001000101110" when 1322,
"1110011101111111" when 1323,
"0001111111111100" when 1324,
"0011111101110011" when 1325,
"0010110101000100" when 1326,
"1111011110101010" when 1327,
"1100100010010110" when 1328,
"1100010011011110" when 1329,
"1110111101101100" when 1330,
"0010011011110010" when 1331,
"0011111111111111" when 1332,
"0010011011111001" when 1333,
"1110111101110100" when 1334,
"1100010011100001" when 1335,
"1100100010010001" when 1336,
"1111011110100010" when 1337,
"0010110100111110" when 1338,
"0011111101110100" when 1339,
"0010000000000011" when 1340,
"1110011110000110" when 1341,
"1100001000110000" when 1342,
"1100110100111000" when 1343,
"1111111111111100" when 1344,
"0011001011000011" when 1345,
"0011110111010010" when 1346,
"0001100010000001" when 1347,
"1110000000000100" when 1348,
"1100000010001101" when 1349,
"1101001010111100" when 1350,
"0000100001010110" when 1351,
"0011011101101010" when 1352,
"0011101100100010" when 1353,
"0001000010010100" when 1354,
"1101100100001110" when 1355,
"1100000000000001" when 1356,
"1101100100000111" when 1357,
"0001000010001100" when 1358,
"0011101100011111" when 1359,
"0011011101101111" when 1360,
"0000100001011110" when 1361,
"1101001011000010" when 1362,
"1100000010001100" when 1363,
"1101111111111101" when 1364,
"0001100001111001" when 1365,
"0011110111010000" when 1366,
"0011001011001000" when 1367,
"0000000000000100" when 1368,
"1100110100111101" when 1369,
"1100001000101110" when 1370,
"1110011101111111" when 1371,
"0001111111111100" when 1372,
"0011111101110011" when 1373,
"0010110101000100" when 1374,
"1111011110101010" when 1375,
"1100100010010110" when 1376,
"1100010011011110" when 1377,
"1110111101101100" when 1378,
"0010011011110010" when 1379,
"0011111111111111" when 1380,
"0010011011111001" when 1381,
"1110111101110100" when 1382,
"1100010011100001" when 1383,
"1100100010010001" when 1384,
"1111011110100010" when 1385,
"0010110100111110" when 1386,
"0011111101110100" when 1387,
"0010000000000011" when 1388,
"1110011110000111" when 1389,
"1100001000110000" when 1390,
"1100110100111000" when 1391,
"1111111111111100" when 1392,
"0011001011000011" when 1393,
"0011110111010010" when 1394,
"0001100010000001" when 1395,
"1110000000000100" when 1396,
"1100000010001101" when 1397,
"1101001010111100" when 1398,
"0000100001010110" when 1399,
"0011011101101010" when 1400,
"0011101100100010" when 1401,
"0001000010010100" when 1402,
"1101100100001110" when 1403,
"1100000000000001" when 1404,
"1101100100000111" when 1405,
"0001000010001100" when 1406,
"0011101100011111" when 1407,
"0011011101101111" when 1408,
"0000100001011110" when 1409,
"1101001011000010" when 1410,
"1100000010001100" when 1411,
"1101111111111101" when 1412,
"0001100001111001" when 1413,
"0011110111010000" when 1414,
"0011001011001000" when 1415,
"0000000000000100" when 1416,
"1100110100111101" when 1417,
"1100001000101110" when 1418,
"1110011101111111" when 1419,
"0001111111111100" when 1420,
"0011111101110011" when 1421,
"0010110101000100" when 1422,
"1111011110101010" when 1423,
"1100100010010110" when 1424,
"1100010011011110" when 1425,
"1110111101101100" when 1426,
"0010011011110010" when 1427,
"0011111111111111" when 1428,
"0010011011111001" when 1429,
"1110111101110100" when 1430,
"1100010011100001" when 1431,
"1100100010010001" when 1432,
"1111011110100010" when 1433,
"0010110100111110" when 1434,
"0011111101110100" when 1435,
"0010000000000011" when 1436,
"1110011110000111" when 1437,
"1100001000110000" when 1438,
"1100110100110111" when 1439,
"1111111111111100" when 1440,
"0011001011000011" when 1441,
"0011110111010010" when 1442,
"0001100010000010" when 1443,
"1110000000000100" when 1444,
"1100000010001101" when 1445,
"1101001010111100" when 1446,
"0000100001010110" when 1447,
"0011011101101010" when 1448,
"0011101100100010" when 1449,
"0001000010010100" when 1450,
"1101100100001110" when 1451,
"1100000000000001" when 1452,
"1101100100000111" when 1453,
"0001000010001100" when 1454,
"0011101100011111" when 1455,
"0011011101101111" when 1456,
"0000100001011111" when 1457,
"1101001011000010" when 1458,
"1100000010001100" when 1459,
"1101111111111101" when 1460,
"0001100001111001" when 1461,
"0011110111010000" when 1462,
"0011001011001001" when 1463,
"0000000000000100" when 1464,
"1100110100111101" when 1465,
"1100001000101110" when 1466,
"1110011101111110" when 1467,
"0001111111111100" when 1468,
"0011111101110011" when 1469,
"0010110101000100" when 1470,
"1111011110101011" when 1471,
"1100100010010110" when 1472,
"1100010011011110" when 1473,
"1110111101101100" when 1474,
"0010011011110010" when 1475,
"0011111111111111" when 1476,
"0010011011111001" when 1477,
"1110111101110100" when 1478,
"1100010011100001" when 1479,
"1100100010010001" when 1480,
"1111011110100001" when 1481,
"0010110100111101" when 1482,
"0011111101110100" when 1483,
"0010000000000100" when 1484,
"1110011110000111" when 1485,
"1100001000110000" when 1486,
"1100110100110111" when 1487,
"1111111111111100" when 1488,
"0011001011000011" when 1489,
"0011110111010010" when 1490,
"0001100010000010" when 1491,
"1110000000000101" when 1492,
"1100000010001101" when 1493,
"1101001010111100" when 1494,
"0000100001010101" when 1495,
"0011011101101010" when 1496,
"0011101100100010" when 1497,
"0001000010010101" when 1498,
"1101100100001110" when 1499,
"1100000000000001" when 1500,
"1101100100000111" when 1501,
"0001000010001011" when 1502,
"0011101100011111" when 1503,
"0011011101101111" when 1504,
"0000100001011111" when 1505,
"1101001011000011" when 1506,
"1100000010001100" when 1507,
"1101111111111100" when 1508,
"0001100001111001" when 1509,
"0011110111010000" when 1510,
"0011001011001001" when 1511,
"0000000000000100" when 1512,
"1100110100111101" when 1513,
"1100001000101110" when 1514,
"1110011101111110" when 1515,
"0001111111111011" when 1516,
"0011111101110011" when 1517,
"0010110101000100" when 1518,
"1111011110101011" when 1519,
"1100100010010110" when 1520,
"1100010011011110" when 1521,
"1110111101101011" when 1522,
"0010011011110010" when 1523,
"0011111111111111" when 1524,
"0010011011111001" when 1525,
"1110111101110101" when 1526,
"1100010011100001" when 1527,
"1100100010010001" when 1528,
"1111011110100001" when 1529,
"0010110100111101" when 1530,
"0011111101110100" when 1531,
"0010000000000100" when 1532,
"1110011110000111" when 1533,
"1100001000110000" when 1534,
"1100110100110111" when 1535,
"1111111111111100" when 1536,
"0011001011000011" when 1537,
"0011110111010010" when 1538,
"0001100010000010" when 1539,
"1110000000000101" when 1540,
"1100000010001101" when 1541,
"1101001010111100" when 1542,
"0000100001010101" when 1543,
"0011011101101010" when 1544,
"0011101100100010" when 1545,
"0001000010010101" when 1546,
"1101100100001110" when 1547,
"1100000000000001" when 1548,
"1101100100000111" when 1549,
"0001000010001011" when 1550,
"0011101100011110" when 1551,
"0011011101101111" when 1552,
"0000100001011111" when 1553,
"1101001011000011" when 1554,
"1100000010001100" when 1555,
"1101111111111100" when 1556,
"0001100001111001" when 1557,
"0011110111010000" when 1558,
"0011001011001001" when 1559,
"0000000000000100" when 1560,
"1100110100111101" when 1561,
"1100001000101110" when 1562,
"1110011101111110" when 1563,
"0001111111111011" when 1564,
"0011111101110011" when 1565,
"0010110101000100" when 1566,
"1111011110101011" when 1567,
"1100100010010110" when 1568,
"1100010011011110" when 1569,
"1110111101101011" when 1570,
"0010011011110010" when 1571,
"0011111111111111" when 1572,
"0010011011111001" when 1573,
"1110111101110101" when 1574,
"1100010011100010" when 1575,
"1100100010010001" when 1576,
"1111011110100001" when 1577,
"0010110100111101" when 1578,
"0011111101110100" when 1579,
"0010000000000100" when 1580,
"1110011110000111" when 1581,
"1100001000110000" when 1582,
"1100110100110111" when 1583,
"1111111111111100" when 1584,
"0011001011000011" when 1585,
"0011110111010011" when 1586,
"0001100010000010" when 1587,
"1110000000000101" when 1588,
"1100000010001101" when 1589,
"1101001010111100" when 1590,
"0000100001010101" when 1591,
"0011011101101010" when 1592,
"0011101100100010" when 1593,
"0001000010010101" when 1594,
"1101100100001111" when 1595,
"1100000000000001" when 1596,
"1101100100000111" when 1597,
"0001000010001011" when 1598,
"0011101100011110" when 1599,
"0011011101101111" when 1600,
"0000100001011111" when 1601,
"1101001011000011" when 1602,
"1100000010001100" when 1603,
"1101111111111100" when 1604,
"0001100001111001" when 1605,
"0011110111010000" when 1606,
"0011001011001001" when 1607,
"0000000000000101" when 1608,
"1100110100111101" when 1609,
"1100001000101101" when 1610,
"1110011101111110" when 1611,
"0001111111111011" when 1612,
"0011111101110011" when 1613,
"0010110101000100" when 1614,
"1111011110101011" when 1615,
"1100100010010110" when 1616,
"1100010011011110" when 1617,
"1110111101101011" when 1618,
"0010011011110001" when 1619,
"0011111111111111" when 1620,
"0010011011111001" when 1621,
"1110111101110101" when 1622,
"1100010011100010" when 1623,
"1100100010010001" when 1624,
"1111011110100001" when 1625,
"0010110100111101" when 1626,
"0011111101110100" when 1627,
"0010000000000100" when 1628,
"1110011110000111" when 1629,
"1100001000110000" when 1630,
"1100110100110111" when 1631,
"1111111111111011" when 1632,
"0011001011000011" when 1633,
"0011110111010011" when 1634,
"0001100010000010" when 1635,
"1110000000000101" when 1636,
"1100000010001101" when 1637,
"1101001010111100" when 1638,
"0000100001010101" when 1639,
"0011011101101010" when 1640,
"0011101100100010" when 1641,
"0001000010010101" when 1642,
"1101100100001111" when 1643,
"1100000000000001" when 1644,
"1101100100000110" when 1645,
"0001000010001011" when 1646,
"0011101100011110" when 1647,
"0011011101101111" when 1648,
"0000100001011111" when 1649,
"1101001011000011" when 1650,
"1100000010001100" when 1651,
"1101111111111100" when 1652,
"0001100001111001" when 1653,
"0011110111010000" when 1654,
"0011001011001001" when 1655,
"0000000000000101" when 1656,
"1100110100111101" when 1657,
"1100001000101101" when 1658,
"1110011101111110" when 1659,
"0001111111111011" when 1660,
"0011111101110011" when 1661,
"0010110101000100" when 1662,
"1111011110101011" when 1663,
"1100100010010110" when 1664,
"1100010011011110" when 1665,
"1110111101101011" when 1666,
"0010011011110001" when 1667,
"0011111111111111" when 1668,
"0010011011111010" when 1669,
"1110111101110101" when 1670,
"1100010011100010" when 1671,
"1100100010010001" when 1672,
"1111011110100001" when 1673,
"0010110100111101" when 1674,
"0011111101110100" when 1675,
"0010000000000100" when 1676,
"1110011110000111" when 1677,
"1100001000110000" when 1678,
"1100110100110111" when 1679,
"1111111111111011" when 1680,
"0011001011000011" when 1681,
"0011110111010011" when 1682,
"0001100010000010" when 1683,
"1110000000000101" when 1684,
"1100000010001101" when 1685,
"1101001010111100" when 1686,
"0000100001010101" when 1687,
"0011011101101010" when 1688,
"0011101100100010" when 1689,
"0001000010010101" when 1690,
"1101100100001111" when 1691,
"1100000000000001" when 1692,
"1101100100000110" when 1693,
"0001000010001011" when 1694,
"0011101100011110" when 1695,
"0011011101101111" when 1696,
"0000100001011111" when 1697,
"1101001011000011" when 1698,
"1100000010001100" when 1699,
"1101111111111100" when 1700,
"0001100001111000" when 1701,
"0011110111010000" when 1702,
"0011001011001001" when 1703,
"0000000000000101" when 1704,
"1100110100111101" when 1705,
"1100001000101101" when 1706,
"1110011101111110" when 1707,
"0001111111111011" when 1708,
"0011111101110011" when 1709,
"0010110101000101" when 1710,
"1111011110101011" when 1711,
"1100100010010110" when 1712,
"1100010011011110" when 1713,
"1110111101101011" when 1714,
"0010011011110001" when 1715,
"0011111111111111" when 1716,
"0010011011111010" when 1717,
"1110111101110101" when 1718,
"1100010011100010" when 1719,
"1100100010010001" when 1720,
"1111011110100001" when 1721,
"0010110100111101" when 1722,
"0011111101110100" when 1723,
"0010000000000100" when 1724,
"1110011110001000" when 1725,
"1100001000110000" when 1726,
"1100110100110111" when 1727,
"1111111111111011" when 1728,
"0011001011000011" when 1729,
"0011110111010011" when 1730,
"0001100010000010" when 1731,
"1110000000000101" when 1732,
"1100000010001101" when 1733,
"1101001010111011" when 1734,
"0000100001010101" when 1735,
"0011011101101010" when 1736,
"0011101100100010" when 1737,
"0001000010010101" when 1738,
"1101100100001111" when 1739,
"1100000000000001" when 1740,
"1101100100000110" when 1741,
"0001000010001011" when 1742,
"0011101100011110" when 1743,
"0011011101101111" when 1744,
"0000100001011111" when 1745,
"1101001011000011" when 1746,
"1100000010001100" when 1747,
"1101111111111100" when 1748,
"0001100001111000" when 1749,
"0011110111010000" when 1750,
"0011001011001001" when 1751,
"0000000000000101" when 1752,
"1100110100111110" when 1753,
"1100001000101101" when 1754,
"1110011101111110" when 1755,
"0001111111111011" when 1756,
"0011111101110011" when 1757,
"0010110101000101" when 1758,
"1111011110101011" when 1759,
"1100100010010110" when 1760,
"1100010011011110" when 1761,
"1110111101101011" when 1762,
"0010011011110001" when 1763,
"0011111111111111" when 1764,
"0010011011111010" when 1765,
"1110111101110101" when 1766,
"1100010011100010" when 1767,
"1100100010010001" when 1768,
"1111011110100000" when 1769,
"0010110100111101" when 1770,
"0011111101110100" when 1771,
"0010000000000100" when 1772,
"1110011110001000" when 1773,
"1100001000110000" when 1774,
"1100110100110111" when 1775,
"1111111111111011" when 1776,
"0011001011000010" when 1777,
"0011110111010011" when 1778,
"0001100010000011" when 1779,
"1110000000000101" when 1780,
"1100000010001101" when 1781,
"1101001010111011" when 1782,
"0000100001010101" when 1783,
"0011011101101010" when 1784,
"0011101100100010" when 1785,
"0001000010010101" when 1786,
"1101100100001111" when 1787,
"1100000000000001" when 1788,
"1101100100000110" when 1789,
"0001000010001011" when 1790,
"0011101100011110" when 1791,
"0011011101101111" when 1792,
"0000100001100000" when 1793,
"1101001011000011" when 1794,
"1100000010001100" when 1795,
"1101111111111100" when 1796,
"0001100001111000" when 1797,
"0011110111010000" when 1798,
"0011001011001001" when 1799,
"0000000000000101" when 1800,
"1100110100111110" when 1801,
"1100001000101101" when 1802,
"1110011101111101" when 1803,
"0001111111111011" when 1804,
"0011111101110011" when 1805,
"0010110101000101" when 1806,
"1111011110101100" when 1807,
"1100100010010110" when 1808,
"1100010011011101" when 1809,
"1110111101101011" when 1810,
"0010011011110001" when 1811,
"0011111111111111" when 1812,
"0010011011111010" when 1813,
"1110111101110101" when 1814,
"1100010011100010" when 1815,
"1100100010010001" when 1816,
"1111011110100000" when 1817,
"0010110100111101" when 1818,
"0011111101110100" when 1819,
"0010000000000100" when 1820,
"1110011110001000" when 1821,
"1100001000110000" when 1822,
"1100110100110111" when 1823,
"1111111111111011" when 1824,
"0011001011000010" when 1825,
"0011110111010011" when 1826,
"0001100010000011" when 1827,
"1110000000000101" when 1828,
"1100000010001101" when 1829,
"1101001010111011" when 1830,
"0000100001010100" when 1831,
"0011011101101010" when 1832,
"0011101100100011" when 1833,
"0001000010010110" when 1834,
"1101100100001111" when 1835,
"1100000000000001" when 1836,
"1101100100000110" when 1837,
"0001000010001010" when 1838,
"0011101100011110" when 1839,
"0011011101101111" when 1840,
"0000100001100000" when 1841,
"1101001011000011" when 1842,
"1100000010001100" when 1843,
"1101111111111100" when 1844,
"0001100001111000" when 1845,
"0011110111010000" when 1846,
"0011001011001001" when 1847,
"0000000000000101" when 1848,
"1100110100111110" when 1849,
"1100001000101101" when 1850,
"1110011101111101" when 1851,
"0001111111111010" when 1852,
"0011111101110011" when 1853,
"0010110101000101" when 1854,
"1111011110101100" when 1855,
"1100100010010110" when 1856,
"1100010011011101" when 1857,
"1110111101101010" when 1858,
"0010011011110001" when 1859,
"0011111111111111" when 1860,
"0010011011111010" when 1861,
"1110111101110110" when 1862,
"1100010011100010" when 1863,
"1100100010010001" when 1864,
"1111011110100000" when 1865,
"0010110100111101" when 1866,
"0011111101110100" when 1867,
"0010000000000101" when 1868,
"1110011110001000" when 1869,
"1100001000110000" when 1870,
"1100110100110111" when 1871,
"1111111111111011" when 1872,
"0011001011000010" when 1873,
"0011110111010011" when 1874,
"0001100010000011" when 1875,
"1110000000000110" when 1876,
"1100000010001101" when 1877,
"1101001010111011" when 1878,
"0000100001010100" when 1879,
"0011011101101010" when 1880,
"0011101100100011" when 1881,
"0001000010010110" when 1882,
"1101100100001111" when 1883,
"1100000000000001" when 1884,
"1101100100000110" when 1885,
"0001000010001010" when 1886,
"0011101100011110" when 1887,
"0011011101101111" when 1888,
"0000100001100000" when 1889,
"1101001011000011" when 1890,
"1100000010001100" when 1891,
"1101111111111011" when 1892,
"0001100001111000" when 1893,
"0011110111010000" when 1894,
"0011001011001001" when 1895,
"0000000000000101" when 1896,
"1100110100111110" when 1897,
"1100001000101101" when 1898,
"1110011101111101" when 1899,
"0001111111111010" when 1900,
"0011111101110011" when 1901,
"0010110101000101" when 1902,
"1111011110101100" when 1903,
"1100100010010111" when 1904,
"1100010011011101" when 1905,
"1110111101101010" when 1906,
"0010011011110001" when 1907,
"0011111111111111" when 1908,
"0010011011111010" when 1909,
"1110111101110110" when 1910,
"1100010011100010" when 1911,
"1100100010010001" when 1912,
"1111011110100000" when 1913,
"0010110100111101" when 1914,
"0011111101110100" when 1915,
"0010000000000101" when 1916,
"1110011110001000" when 1917,
"1100001000110000" when 1918,
"1100110100110111" when 1919,
"1111111111111011" when 1920,
"0011001011000010" when 1921,
"0011110111010011" when 1922,
"0001100010000011" when 1923,
"1110000000000110" when 1924,
"1100000010001101" when 1925,
"1101001010111011" when 1926,
"0000100001010100" when 1927,
"0011011101101001" when 1928,
"0011101100100011" when 1929,
"0001000010010110" when 1930,
"1101100100001111" when 1931,
"1100000000000001" when 1932,
"1101100100000110" when 1933,
"0001000010001010" when 1934,
"0011101100011110" when 1935,
"0011011101101111" when 1936,
"0000100001100000" when 1937,
"1101001011000100" when 1938,
"1100000010001100" when 1939,
"1101111111111011" when 1940,
"0001100001111000" when 1941,
"0011110111010000" when 1942,
"0011001011001001" when 1943,
"0000000000000110" when 1944,
"1100110100111110" when 1945,
"1100001000101101" when 1946,
"1110011101111101" when 1947,
"0001111111111010" when 1948,
"0011111101110011" when 1949,
"0010110101000101" when 1950,
"1111011110101100" when 1951,
"1100100010010111" when 1952,
"1100010011011101" when 1953,
"1110111101101010" when 1954,
"0010011011110001" when 1955,
"0011111111111111" when 1956,
"0010011011111010" when 1957,
"1110111101110110" when 1958,
"1100010011100010" when 1959,
"1100100010010000" when 1960,
"1111011110100000" when 1961,
"0010110100111100" when 1962,
"0011111101110100" when 1963,
"0010000000000101" when 1964,
"1110011110001000" when 1965,
"1100001000110000" when 1966,
"1100110100110110" when 1967,
"1111111111111010" when 1968,
"0011001011000010" when 1969,
"0011110111010011" when 1970,
"0001100010000011" when 1971,
"1110000000000110" when 1972,
"1100000010001101" when 1973,
"1101001010111011" when 1974,
"0000100001010100" when 1975,
"0011011101101001" when 1976,
"0011101100100011" when 1977,
"0001000010010110" when 1978,
"1101100100001111" when 1979,
"1100000000000001" when 1980,
"1101100100000110" when 1981,
"0001000010001010" when 1982,
"0011101100011110" when 1983,
"0011011101110000" when 1984,
"0000100001100000" when 1985,
"1101001011000100" when 1986,
"1100000010001100" when 1987,
"1101111111111011" when 1988,
"0001100001111000" when 1989,
"0011110111010000" when 1990,
"0011001011001010" when 1991,
"0000000000000110" when 1992,
"1100110100111110" when 1993,
"1100001000101101" when 1994,
"1110011101111101" when 1995,
"0001111111111010" when 1996,
"0011111101110011" when 1997,
"0010110101000101" when 1998,
"1111011110101100" when 1999,
"1100100010010111" when 2000,
"1100010011011101" when 2001,
"1110111101101010" when 2002,
"0010011011110000" when 2003,
"0011111111111111" when 2004,
"0010011011111010" when 2005,
"1110111101110110" when 2006,
"1100010011100010" when 2007,
"1100100010010000" when 2008,
"1111011110100000" when 2009,
"0010110100111100" when 2010,
"0011111101110100" when 2011,
"0010000000000101" when 2012,
"1110011110001000" when 2013,
"1100001000110000" when 2014,
"1100110100110110" when 2015,
"1111111111111010" when 2016,
"0011001011000010" when 2017,
"0011110111010011" when 2018,
"0001100010000011" when 2019,
"1110000000000110" when 2020,
"1100000010001101" when 2021,
"1101001010111011" when 2022,
"0000100001010100" when 2023,
"0011011101101001" when 2024,
"0011101100100011" when 2025,
"0001000010010110" when 2026,
"1101100100010000" when 2027,
"1100000000000001" when 2028,
"1101100100000110" when 2029,
"0001000010001010" when 2030,
"0011101100011110" when 2031,
"0011011101110000" when 2032,
"0000100001100000" when 2033,
"1101001011000100" when 2034,
"1100000010001100" when 2035,
"1101111111111011" when 2036,
"0001100001111000" when 2037,
"0011110111010000" when 2038,
"0011001011001010" when 2039,
"0000000000000110" when 2040,
"1100110100111110" when 2041,
"1100001000101101" when 2042,
"1110011101111101" when 2043,
"0001111111111010" when 2044,
"0011111101110010" when 2045,
"0010110101000101" when 2046,
"1111011110101100" when 2047,
"1100100010010111" when 2048,
"1100010011011101" when 2049,
"1110111101101010" when 2050,
"0010011011110000" when 2051,
"0011111111111111" when 2052,
"0010011011111011" when 2053,
"1110111101110110" when 2054,
"1100010011100010" when 2055,
"1100100010010000" when 2056,
"1111011110100000" when 2057,
"0010110100111100" when 2058,
"0011111101110100" when 2059,
"0010000000000101" when 2060,
"1110011110001001" when 2061,
"1100001000110000" when 2062,
"1100110100110110" when 2063,
"1111111111111010" when 2064,
"0011001011000010" when 2065,
"0011110111010011" when 2066,
"0001100010000011" when 2067,
"1110000000000110" when 2068,
"1100000010001110" when 2069,
"1101001010111011" when 2070,
"0000100001010100" when 2071,
"0011011101101001" when 2072,
"0011101100100011" when 2073,
"0001000010010110" when 2074,
"1101100100010000" when 2075,
"1100000000000001" when 2076,
"1101100100000101" when 2077,
"0001000010001010" when 2078,
"0011101100011110" when 2079,
"0011011101110000" when 2080,
"0000100001100000" when 2081,
"1101001011000100" when 2082,
"1100000010001100" when 2083,
"1101111111111011" when 2084,
"0001100001110111" when 2085,
"0011110111010000" when 2086,
"0011001011001010" when 2087,
"0000000000000110" when 2088,
"1100110100111110" when 2089,
"1100001000101101" when 2090,
"1110011101111101" when 2091,
"0001111111111010" when 2092,
"0011111101110010" when 2093,
"0010110101000101" when 2094,
"1111011110101100" when 2095,
"1100100010010111" when 2096,
"1100010011011101" when 2097,
"1110111101101010" when 2098,
"0010011011110000" when 2099,
"0011111111111111" when 2100,
"0010011011111011" when 2101,
"1110111101110110" when 2102,
"1100010011100010" when 2103,
"1100100010010000" when 2104,
"1111011110011111" when 2105,
"0010110100111100" when 2106,
"0011111101110100" when 2107,
"0010000000000101" when 2108,
"1110011110001001" when 2109,
"1100001000110000" when 2110,
"1100110100110110" when 2111,
"1111111111111010" when 2112,
"0011001011000010" when 2113,
"0011110111010011" when 2114,
"0001100010000011" when 2115,
"1110000000000110" when 2116,
"1100000010001110" when 2117,
"1101001010111011" when 2118,
"0000100001010011" when 2119,
"0011011101101001" when 2120,
"0011101100100011" when 2121,
"0001000010010110" when 2122,
"1101100100010000" when 2123,
"1100000000000001" when 2124,
"1101100100000101" when 2125,
"0001000010001010" when 2126,
"0011101100011110" when 2127,
"0011011101110000" when 2128,
"0000100001100001" when 2129,
"1101001011000100" when 2130,
"1100000010001100" when 2131,
"1101111111111011" when 2132,
"0001100001110111" when 2133,
"0011110111010000" when 2134,
"0011001011001010" when 2135,
"0000000000000110" when 2136,
"1100110100111110" when 2137,
"1100001000101101" when 2138,
"1110011101111100" when 2139,
"0001111111111010" when 2140,
"0011111101110010" when 2141,
"0010110101000101" when 2142,
"1111011110101101" when 2143,
"1100100010010111" when 2144,
"1100010011011101" when 2145,
"1110111101101010" when 2146,
"0010011011110000" when 2147,
"0011111111111111" when 2148,
"0010011011111011" when 2149,
"1110111101110110" when 2150,
"1100010011100010" when 2151,
"1100100010010000" when 2152,
"1111011110011111" when 2153,
"0010110100111100" when 2154,
"0011111101110100" when 2155,
"0010000000000101" when 2156,
"1110011110001001" when 2157,
"1100001000110001" when 2158,
"1100110100110110" when 2159,
"1111111111111010" when 2160,
"0011001011000010" when 2161,
"0011110111010011" when 2162,
"0001100010000100" when 2163,
"1110000000000110" when 2164,
"1100000010001110" when 2165,
"1101001010111010" when 2166,
"0000100001010011" when 2167,
"0011011101101001" when 2168,
"0011101100100011" when 2169,
"0001000010010111" when 2170,
"1101100100010000" when 2171,
"1100000000000001" when 2172,
"1101100100000101" when 2173,
"0001000010001001" when 2174,
"0011101100011110" when 2175,
"0011011101110000" when 2176,
"0000100001100001" when 2177,
"1101001011000100" when 2178,
"1100000010001100" when 2179,
"1101111111111011" when 2180,
"0001100001110111" when 2181,
"0011110111001111" when 2182,
"0011001011001010" when 2183,
"0000000000000110" when 2184,
"1100110100111110" when 2185,
"1100001000101101" when 2186,
"1110011101111100" when 2187,
"0001111111111010" when 2188,
"0011111101110010" when 2189,
"0010110101000110" when 2190,
"1111011110101101" when 2191,
"1100100010010111" when 2192,
"1100010011011101" when 2193,
"1110111101101001" when 2194,
"0010011011110000" when 2195,
"0011111111111111" when 2196,
"0010011011111011" when 2197,
"1110111101110111" when 2198,
"1100010011100010" when 2199,
"1100100010010000" when 2200,
"1111011110011111" when 2201,
"0010110100111100" when 2202,
"0011111101110100" when 2203,
"0010000000000101" when 2204,
"1110011110001001" when 2205,
"1100001000110001" when 2206,
"1100110100110110" when 2207,
"1111111111111010" when 2208,
"0011001011000010" when 2209,
"0011110111010011" when 2210,
"0001100010000100" when 2211,
"1110000000000110" when 2212,
"1100000010001110" when 2213,
"1101001010111010" when 2214,
"0000100001010011" when 2215,
"0011011101101001" when 2216,
"0011101100100011" when 2217,
"0001000010010111" when 2218,
"1101100100010000" when 2219,
"1100000000000001" when 2220,
"1101100100000101" when 2221,
"0001000010001001" when 2222,
"0011101100011110" when 2223,
"0011011101110000" when 2224,
"0000100001100001" when 2225,
"1101001011000100" when 2226,
"1100000010001100" when 2227,
"1101111111111010" when 2228,
"0001100001110111" when 2229,
"0011110111001111" when 2230,
"0011001011001010" when 2231,
"0000000000000110" when 2232,
"1100110100111110" when 2233,
"1100001000101101" when 2234,
"1110011101111100" when 2235,
"0001111111111001" when 2236,
"0011111101110010" when 2237,
"0010110101000110" when 2238,
"1111011110101101" when 2239,
"1100100010010111" when 2240,
"1100010011011101" when 2241,
"1110111101101001" when 2242,
"0010011011110000" when 2243,
"0011111111111111" when 2244,
"0010011011111011" when 2245,
"1110111101110111" when 2246,
"1100010011100010" when 2247,
"1100100010010000" when 2248,
"1111011110011111" when 2249,
"0010110100111100" when 2250,
"0011111101110100" when 2251,
"0010000000000110" when 2252,
"1110011110001001" when 2253,
"1100001000110001" when 2254,
"1100110100110110" when 2255,
"1111111111111001" when 2256,
"0011001011000010" when 2257,
"0011110111010011" when 2258,
"0001100010000100" when 2259,
"1110000000000111" when 2260,
"1100000010001110" when 2261,
"1101001010111010" when 2262,
"0000100001010011" when 2263,
"0011011101101001" when 2264,
"0011101100100011" when 2265,
"0001000010010111" when 2266,
"1101100100010000" when 2267,
"1100000000000001" when 2268,
"1101100100000101" when 2269,
"0001000010001001" when 2270,
"0011101100011110" when 2271,
"0011011101110000" when 2272,
"0000100001100001" when 2273,
"1101001011000100" when 2274,
"1100000010001100" when 2275,
"1101111111111010" when 2276,
"0001100001110111" when 2277,
"0011110111001111" when 2278,
"0011001011001010" when 2279,
"0000000000000111" when 2280,
"1100110100111111" when 2281,
"1100001000101101" when 2282,
"1110011101111100" when 2283,
"0001111111111001" when 2284,
"0011111101110010" when 2285,
"0010110101000110" when 2286,
"1111011110101101" when 2287,
"1100100010010111" when 2288,
"1100010011011101" when 2289,
"1110111101101001" when 2290,
"0010011011110000" when 2291,
"0011111111111111" when 2292,
"0010011011111011" when 2293,
"1110111101110111" when 2294,
"1100010011100010" when 2295,
"1100100010010000" when 2296,
"1111011110011111" when 2297,
"0010110100111100" when 2298,
"0011111101110100" when 2299,
"0010000000000110" when 2300,
"1110011110001001" when 2301,
"1100001000110001" when 2302,
"1100110100110110" when 2303,
"1111111111111001" when 2304,
"0011001011000001" when 2305,
"0011110111010011" when 2306,
"0001100010000100" when 2307,
"1110000000000111" when 2308,
"1100000010001110" when 2309,
"1101001010111010" when 2310,
"0000100001010011" when 2311,
"0011011101101001" when 2312,
"0011101100100011" when 2313,
"0001000010010111" when 2314,
"1101100100010000" when 2315,
"1100000000000001" when 2316,
"1101100100000101" when 2317,
"0001000010001001" when 2318,
"0011101100011110" when 2319,
"0011011101110000" when 2320,
"0000100001100001" when 2321,
"1101001011000100" when 2322,
"1100000010001100" when 2323,
"1101111111111010" when 2324,
"0001100001110111" when 2325,
"0011110111001111" when 2326,
"0011001011001010" when 2327,
"0000000000000111" when 2328,
"1100110100111111" when 2329,
"1100001000101101" when 2330,
"1110011101111100" when 2331,
"0001111111111001" when 2332,
"0011111101110010" when 2333,
"0010110101000110" when 2334,
"1111011110101101" when 2335,
"1100100010010111" when 2336,
"1100010011011101" when 2337,
"1110111101101001" when 2338,
"0010011011110000" when 2339,
"0011111111111111" when 2340,
"0010011011111011" when 2341,
"1110111101110111" when 2342,
"1100010011100010" when 2343,
"1100100010010000" when 2344,
"1111011110011111" when 2345,
"0010110100111100" when 2346,
"0011111101110100" when 2347,
"0010000000000110" when 2348,
"1110011110001001" when 2349,
"1100001000110001" when 2350,
"1100110100110110" when 2351,
"1111111111111001" when 2352,
"0011001011000001" when 2353,
"0011110111010011" when 2354,
"0001100010000100" when 2355,
"1110000000000111" when 2356,
"1100000010001110" when 2357,
"1101001010111010" when 2358,
"0000100001010011" when 2359,
"0011011101101001" when 2360,
"0011101100100011" when 2361,
"0001000010010111" when 2362,
"1101100100010000" when 2363,
"1100000000000001" when 2364,
"1101100100000101" when 2365,
"0001000010001001" when 2366,
"0011101100011110" when 2367,
"0011011101110000" when 2368,
"0000100001100001" when 2369,
"1101001011000100" when 2370,
"1100000010001100" when 2371,
"1101111111111010" when 2372,
"0001100001110111" when 2373,
"0011110111001111" when 2374,
"0011001011001010" when 2375,
"0000000000000111" when 2376,
"1100110100111111" when 2377,
"1100001000101101" when 2378,
"1110011101111100" when 2379,
"0001111111111001" when 2380,
"0011111101110010" when 2381,
"0010110101000110" when 2382,
"1111011110101101" when 2383,
"1100100010010111" when 2384,
"1100010011011101" when 2385,
"1110111101101001" when 2386,
"0010011011110000" when 2387,
"0011111111111111" when 2388,
"0010011011111011" when 2389,
"1110111101110111" when 2390,
"1100010011100011" when 2391,
"1100100010010000" when 2392,
"1111011110011111" when 2393,
"0010110100111011" when 2394,
"0011111101110100" when 2395,
"0010000000000110" when 2396,
"1110011110001010" when 2397,
"1100001000110001" when 2398,
"1100110100110110" when 2399,
"1111111111111001" when 2400,
"0011001011000001" when 2401,
"0011110111010011" when 2402,
"0001100010000100" when 2403,
"1110000000000111" when 2404,
"1100000010001110" when 2405,
"1101001010111010" when 2406,
"0000100001010011" when 2407,
"0011011101101001" when 2408,
"0011101100100011" when 2409,
"0001000010010111" when 2410,
"1101100100010001" when 2411,
"1100000000000001" when 2412,
"1101100100000101" when 2413,
"0001000010001001" when 2414,
"0011101100011101" when 2415,
"0011011101110000" when 2416,
"0000100001100010" when 2417,
"1101001011000101" when 2418,
"1100000010001100" when 2419,
"1101111111111010" when 2420,
"0001100001110110" when 2421,
"0011110111001111" when 2422,
"0011001011001010" when 2423,
"0000000000000111" when 2424,
"1100110100111111" when 2425,
"1100001000101101" when 2426,
"1110011101111100" when 2427,
"0001111111111001" when 2428,
"0011111101110010" when 2429,
"0010110101000110" when 2430,
"1111011110101101" when 2431,
"1100100010010111" when 2432,
"1100010011011101" when 2433,
"1110111101101001" when 2434,
"0010011011101111" when 2435,
"0011111111111111" when 2436,
"0010011011111011" when 2437,
"1110111101110111" when 2438,
"1100010011100011" when 2439,
"1100100010010000" when 2440,
"1111011110011110" when 2441,
"0010110100111011" when 2442,
"0011111101110100" when 2443,
"0010000000000110" when 2444,
"1110011110001010" when 2445,
"1100001000110001" when 2446,
"1100110100110110" when 2447,
"1111111111111001" when 2448,
"0011001011000001" when 2449,
"0011110111010011" when 2450,
"0001100010000100" when 2451,
"1110000000000111" when 2452,
"1100000010001110" when 2453,
"1101001010111010" when 2454,
"0000100001010010" when 2455,
"0011011101101001" when 2456,
"0011101100100011" when 2457,
"0001000010010111" when 2458,
"1101100100010001" when 2459,
"1100000000000001" when 2460,
"1101100100000100" when 2461,
"0001000010001001" when 2462,
"0011101100011101" when 2463,
"0011011101110000" when 2464,
"0000100001100010" when 2465,
"1101001011000101" when 2466,
"1100000010001100" when 2467,
"1101111111111010" when 2468,
"0001100001110110" when 2469,
"0011110111001111" when 2470,
"0011001011001010" when 2471,
"0000000000000111" when 2472,
"1100110100111111" when 2473,
"1100001000101101" when 2474,
"1110011101111011" when 2475,
"0001111111111001" when 2476,
"0011111101110010" when 2477,
"0010110101000110" when 2478,
"1111011110101110" when 2479,
"1100100010010111" when 2480,
"1100010011011101" when 2481,
"1110111101101001" when 2482,
"0010011011101111" when 2483,
"0011111111111111" when 2484,
"0010011011111100" when 2485,
"1110111101111000" when 2486,
"1100010011100011" when 2487,
"1100100010010000" when 2488,
"1111011110011110" when 2489,
"0010110100111011" when 2490,
"0011111101110100" when 2491,
"0010000000000110" when 2492,
"1110011110001010" when 2493,
"1100001000110001" when 2494,
"1100110100110101" when 2495,
"1111111111111001" when 2496,
"0011001011000001" when 2497,
"0011110111010011" when 2498,
"0001100010000101" when 2499,
"1110000000000111" when 2500,
"1100000010001110" when 2501,
"1101001010111010" when 2502,
"0000100001010010" when 2503,
"0011011101101001" when 2504,
"0011101100100011" when 2505,
"0001000010011000" when 2506,
"1101100100010001" when 2507,
"1100000000000001" when 2508,
"1101100100000100" when 2509,
"0001000010001000" when 2510,
"0011101100011101" when 2511,
"0011011101110000" when 2512,
"0000100001100010" when 2513,
"1101001011000101" when 2514,
"1100000010001100" when 2515,
"1101111111111010" when 2516,
"0001100001110110" when 2517,
"0011110111001111" when 2518,
"0011001011001011" when 2519,
"0000000000000111" when 2520,
"1100110100111111" when 2521,
"1100001000101101" when 2522,
"1110011101111011" when 2523,
"0001111111111001" when 2524,
"0011111101110010" when 2525,
"0010110101000110" when 2526,
"1111011110101110" when 2527,
"1100100010010111" when 2528,
"1100010011011101" when 2529,
"1110111101101000" when 2530,
"0010011011101111" when 2531,
"0011111111111111" when 2532,
"0010011011111100" when 2533,
"1110111101111000" when 2534,
"1100010011100011" when 2535,
"1100100010010000" when 2536,
"1111011110011110" when 2537,
"0010110100111011" when 2538,
"0011111101110100" when 2539,
"0010000000000110" when 2540,
"1110011110001010" when 2541,
"1100001000110001" when 2542,
"1100110100110101" when 2543,
"1111111111111001" when 2544,
"0011001011000001" when 2545,
"0011110111010011" when 2546,
"0001100010000101" when 2547,
"1110000000000111" when 2548,
"1100000010001110" when 2549,
"1101001010111010" when 2550,
"0000100001010010" when 2551,
"0011011101101000" when 2552,
"0011101100100011" when 2553,
"0001000010011000" when 2554,
"1101100100010001" when 2555,
"1100000000000001" when 2556,
"1101100100000100" when 2557,
"0001000010001000" when 2558,
"0011101100011101" when 2559,
"0011011101110000" when 2560,
"0000100001100010" when 2561,
"1101001011000101" when 2562,
"1100000010001100" when 2563,
"1101111111111010" when 2564,
"0001100001110110" when 2565,
"0011110111001111" when 2566,
"0011001011001011" when 2567,
"0000000000001000" when 2568,
"1100110100111111" when 2569,
"1100001000101101" when 2570,
"1110011101111011" when 2571,
"0001111111111001" when 2572,
"0011111101110010" when 2573,
"0010110101000110" when 2574,
"1111011110101110" when 2575,
"1100100010011000" when 2576,
"1100010011011101" when 2577,
"1110111101101000" when 2578,
"0010011011101111" when 2579,
"0011111111111111" when 2580,
"0010011011111100" when 2581,
"1110111101111000" when 2582,
"1100010011100011" when 2583,
"1100100010010000" when 2584,
"1111011110011110" when 2585,
"0010110100111011" when 2586,
"0011111101110100" when 2587,
"0010000000000110" when 2588,
"1110011110001010" when 2589,
"1100001000110001" when 2590,
"1100110100110101" when 2591,
"1111111111111000" when 2592,
"0011001011000001" when 2593,
"0011110111010011" when 2594,
"0001100010000101" when 2595,
"1110000000001000" when 2596,
"1100000010001110" when 2597,
"1101001010111010" when 2598,
"0000100001010010" when 2599,
"0011011101101000" when 2600,
"0011101100100011" when 2601,
"0001000010011000" when 2602,
"1101100100010001" when 2603,
"1100000000000001" when 2604,
"1101100100000100" when 2605,
"0001000010001000" when 2606,
"0011101100011101" when 2607,
"0011011101110001" when 2608,
"0000100001100010" when 2609,
"1101001011000101" when 2610,
"1100000010001100" when 2611,
"1101111111111001" when 2612,
"0001100001110110" when 2613,
"0011110111001111" when 2614,
"0011001011001011" when 2615,
"0000000000001000" when 2616,
"1100110100111111" when 2617,
"1100001000101101" when 2618,
"1110011101111011" when 2619,
"0001111111111000" when 2620,
"0011111101110010" when 2621,
"0010110101000111" when 2622,
"1111011110101110" when 2623,
"1100100010011000" when 2624,
"1100010011011101" when 2625,
"1110111101101000" when 2626,
"0010011011101111" when 2627,
"0011111111111111" when 2628,
"0010011011111100" when 2629,
"1110111101111000" when 2630,
"1100010011100011" when 2631,
"1100100010001111" when 2632,
"1111011110011110" when 2633,
"0010110100111011" when 2634,
"0011111101110100" when 2635,
"0010000000000111" when 2636,
"1110011110001010" when 2637,
"1100001000110001" when 2638,
"1100110100110101" when 2639,
"1111111111111000" when 2640,
"0011001011000001" when 2641,
"0011110111010011" when 2642,
"0001100010000101" when 2643,
"1110000000001000" when 2644,
"1100000010001110" when 2645,
"1101001010111001" when 2646,
"0000100001010010" when 2647,
"0011011101101000" when 2648,
"0011101100100100" when 2649,
"0001000010011000" when 2650,
"1101100100010001" when 2651,
"1100000000000001" when 2652,
"1101100100000100" when 2653,
"0001000010001000" when 2654,
"0011101100011101" when 2655,
"0011011101110001" when 2656,
"0000100001100010" when 2657,
"1101001011000101" when 2658,
"1100000010001100" when 2659,
"1101111111111001" when 2660,
"0001100001110110" when 2661,
"0011110111001111" when 2662,
"0011001011001011" when 2663,
"0000000000001000" when 2664,
"1100110100111111" when 2665,
"1100001000101101" when 2666,
"1110011101111011" when 2667,
"0001111111111000" when 2668,
"0011111101110010" when 2669,
"0010110101000111" when 2670,
"1111011110101110" when 2671,
"1100100010011000" when 2672,
"1100010011011100" when 2673,
"1110111101101000" when 2674,
"0010011011101111" when 2675,
"0011111111111111" when 2676,
"0010011011111100" when 2677,
"1110111101111000" when 2678,
"1100010011100011" when 2679,
"1100100010001111" when 2680,
"1111011110011110" when 2681,
"0010110100111011" when 2682,
"0011111101110100" when 2683,
"0010000000000111" when 2684,
"1110011110001010" when 2685,
"1100001000110001" when 2686,
"1100110100110101" when 2687,
"1111111111111000" when 2688,
"0011001011000001" when 2689,
"0011110111010011" when 2690,
"0001100010000101" when 2691,
"1110000000001000" when 2692,
"1100000010001110" when 2693,
"1101001010111001" when 2694,
"0000100001010010" when 2695,
"0011011101101000" when 2696,
"0011101100100100" when 2697,
"0001000010011000" when 2698,
"1101100100010001" when 2699,
"1100000000000001" when 2700,
"1101100100000100" when 2701,
"0001000010001000" when 2702,
"0011101100011101" when 2703,
"0011011101110001" when 2704,
"0000100001100010" when 2705,
"1101001011000101" when 2706,
"1100000010001100" when 2707,
"1101111111111001" when 2708,
"0001100001110110" when 2709,
"0011110111001111" when 2710,
"0011001011001011" when 2711,
"0000000000001000" when 2712,
"1100110100111111" when 2713,
"1100001000101101" when 2714,
"1110011101111011" when 2715,
"0001111111111000" when 2716,
"0011111101110010" when 2717,
"0010110101000111" when 2718,
"1111011110101110" when 2719,
"1100100010011000" when 2720,
"1100010011011100" when 2721,
"1110111101101000" when 2722,
"0010011011101111" when 2723,
"0011111111111111" when 2724,
"0010011011111100" when 2725,
"1110111101111000" when 2726,
"1100010011100011" when 2727,
"1100100010001111" when 2728,
"1111011110011110" when 2729,
"0010110100111011" when 2730,
"0011111101110100" when 2731,
"0010000000000111" when 2732,
"1110011110001011" when 2733,
"1100001000110001" when 2734,
"1100110100110101" when 2735,
"1111111111111000" when 2736,
"0011001011000001" when 2737,
"0011110111010011" when 2738,
"0001100010000101" when 2739,
"1110000000001000" when 2740,
"1100000010001110" when 2741,
"1101001010111001" when 2742,
"0000100001010010" when 2743,
"0011011101101000" when 2744,
"0011101100100100" when 2745,
"0001000010011000" when 2746,
"1101100100010001" when 2747,
"1100000000000001" when 2748,
"1101100100000100" when 2749,
"0001000010001000" when 2750,
"0011101100011101" when 2751,
"0011011101110001" when 2752,
"0000100001100011" when 2753,
"1101001011000101" when 2754,
"1100000010001100" when 2755,
"1101111111111001" when 2756,
"0001100001110101" when 2757,
"0011110111001111" when 2758,
"0011001011001011" when 2759,
"0000000000001000" when 2760,
"1100110100111111" when 2761,
"1100001000101101" when 2762,
"1110011101111011" when 2763,
"0001111111111000" when 2764,
"0011111101110010" when 2765,
"0010110101000111" when 2766,
"1111011110101111" when 2767,
"1100100010011000" when 2768,
"1100010011011100" when 2769,
"1110111101101000" when 2770,
"0010011011101111" when 2771,
"0011111111111111" when 2772,
"0010011011111100" when 2773,
"1110111101111000" when 2774,
"1100010011100011" when 2775,
"1100100010001111" when 2776,
"1111011110011101" when 2777,
"0010110100111011" when 2778,
"0011111101110100" when 2779,
"0010000000000111" when 2780,
"1110011110001011" when 2781,
"1100001000110001" when 2782,
"1100110100110101" when 2783,
"1111111111111000" when 2784,
"0011001011000001" when 2785,
"0011110111010011" when 2786,
"0001100010000101" when 2787,
"1110000000001000" when 2788,
"1100000010001110" when 2789,
"1101001010111001" when 2790,
"0000100001010001" when 2791,
"0011011101101000" when 2792,
"0011101100100100" when 2793,
"0001000010011000" when 2794,
"1101100100010001" when 2795,
"1100000000000001" when 2796,
"1101100100000100" when 2797,
"0001000010001000" when 2798,
"0011101100011101" when 2799,
"0011011101110001" when 2800,
"0000100001100011" when 2801,
"1101001011000101" when 2802,
"1100000010001100" when 2803,
"1101111111111001" when 2804,
"0001100001110101" when 2805,
"0011110111001111" when 2806,
"0011001011001011" when 2807,
"0000000000001000" when 2808,
"1100110101000000" when 2809,
"1100001000101101" when 2810,
"1110011101111011" when 2811,
"0001111111111000" when 2812,
"0011111101110010" when 2813,
"0010110101000111" when 2814,
"1111011110101111" when 2815,
"1100100010011000" when 2816,
"1100010011011100" when 2817,
"1110111101101000" when 2818,
"0010011011101110" when 2819,
"0011111111111111" when 2820,
"0010011011111100" when 2821,
"1110111101111001" when 2822,
"1100010011100011" when 2823,
"1100100010001111" when 2824,
"1111011110011101" when 2825,
"0010110100111010" when 2826,
"0011111101110100" when 2827,
"0010000000000111" when 2828,
"1110011110001011" when 2829,
"1100001000110001" when 2830,
"1100110100110101" when 2831,
"1111111111111000" when 2832,
"0011001011000000" when 2833,
"0011110111010100" when 2834,
"0001100010000110" when 2835,
"1110000000001000" when 2836,
"1100000010001110" when 2837,
"1101001010111001" when 2838,
"0000100001010001" when 2839,
"0011011101101000" when 2840,
"0011101100100100" when 2841,
"0001000010011001" when 2842,
"1101100100010010" when 2843,
"1100000000000001" when 2844,
"1101100100000100" when 2845,
"0001000010000111" when 2846,
"0011101100011101" when 2847,
"0011011101110001" when 2848,
"0000100001100011" when 2849,
"1101001011000110" when 2850,
"1100000010001100" when 2851,
"1101111111111001" when 2852,
"0001100001110101" when 2853,
"0011110111001111" when 2854,
"0011001011001011" when 2855,
"0000000000001000" when 2856,
"1100110101000000" when 2857,
"1100001000101100" when 2858,
"1110011101111010" when 2859,
"0001111111111000" when 2860,
"0011111101110010" when 2861,
"0010110101000111" when 2862,
"1111011110101111" when 2863,
"1100100010011000" when 2864,
"1100010011011100" when 2865,
"1110111101100111" when 2866,
"0010011011101110" when 2867,
"0011111111111111" when 2868,
"0010011011111101" when 2869,
"1110111101111001" when 2870,
"1100010011100011" when 2871,
"1100100010001111" when 2872,
"1111011110011101" when 2873,
"0010110100111010" when 2874,
"0011111101110101" when 2875,
"0010000000000111" when 2876,
"1110011110001011" when 2877,
"1100001000110001" when 2878,
"1100110100110101" when 2879,
"1111111111111000" when 2880,
"0011001011000000" when 2881,
"0011110111010100" when 2882,
"0001100010000110" when 2883,
"1110000000001000" when 2884,
"1100000010001110" when 2885,
"1101001010111001" when 2886,
"0000100001010001" when 2887,
"0011011101101000" when 2888,
"0011101100100100" when 2889,
"0001000010011001" when 2890,
"1101100100010010" when 2891,
"1100000000000001" when 2892,
"1101100100000011" when 2893,
"0001000010000111" when 2894,
"0011101100011101" when 2895,
"0011011101110001" when 2896,
"0000100001100011" when 2897,
"1101001011000110" when 2898,
"1100000010001011" when 2899,
"1101111111111001" when 2900,
"0001100001110101" when 2901,
"0011110111001111" when 2902,
"0011001011001011" when 2903,
"0000000000001001" when 2904,
"1100110101000000" when 2905,
"1100001000101100" when 2906,
"1110011101111010" when 2907,
"0001111111111000" when 2908,
"0011111101110010" when 2909,
"0010110101000111" when 2910,
"1111011110101111" when 2911,
"1100100010011000" when 2912,
"1100010011011100" when 2913,
"1110111101100111" when 2914,
"0010011011101110" when 2915,
"0011111111111111" when 2916,
"0010011011111101" when 2917,
"1110111101111001" when 2918,
"1100010011100011" when 2919,
"1100100010001111" when 2920,
"1111011110011101" when 2921,
"0010110100111010" when 2922,
"0011111101110101" when 2923,
"0010000000000111" when 2924,
"1110011110001011" when 2925,
"1100001000110001" when 2926,
"1100110100110101" when 2927,
"1111111111110111" when 2928,
"0011001011000000" when 2929,
"0011110111010100" when 2930,
"0001100010000110" when 2931,
"1110000000001000" when 2932,
"1100000010001110" when 2933,
"1101001010111001" when 2934,
"0000100001010001" when 2935,
"0011011101101000" when 2936,
"0011101100100100" when 2937,
"0001000010011001" when 2938,
"1101100100010010" when 2939,
"1100000000000001" when 2940,
"1101100100000011" when 2941,
"0001000010000111" when 2942,
"0011101100011101" when 2943,
"0011011101110001" when 2944,
"0000100001100011" when 2945,
"1101001011000110" when 2946,
"1100000010001011" when 2947,
"1101111111111001" when 2948,
"0001100001110101" when 2949,
"0011110111001111" when 2950,
"0011001011001011" when 2951,
"0000000000001001" when 2952,
"1100110101000000" when 2953,
"1100001000101100" when 2954,
"1110011101111010" when 2955,
"0001111111111000" when 2956,
"0011111101110010" when 2957,
"0010110101000111" when 2958,
"1111011110101111" when 2959,
"1100100010011000" when 2960,
"1100010011011100" when 2961,
"1110111101100111" when 2962,
"0010011011101110" when 2963,
"0011111111111111" when 2964,
"0010011011111101" when 2965,
"1110111101111001" when 2966,
"1100010011100011" when 2967,
"1100100010001111" when 2968,
"1111011110011101" when 2969,
"0010110100111010" when 2970,
"0011111101110101" when 2971,
"0010000000001000" when 2972,
"1110011110001011" when 2973,
"1100001000110001" when 2974,
"1100110100110101" when 2975,
"1111111111110111" when 2976,
"0011001011000000" when 2977,
"0011110111010100" when 2978,
"0001100010000110" when 2979,
"1110000000001001" when 2980,
"1100000010001110" when 2981,
"1101001010111001" when 2982,
"0000100001010001" when 2983,
"0011011101101000" when 2984,
"0011101100100100" when 2985,
"0001000010011001" when 2986,
"1101100100010010" when 2987,
"1100000000000001" when 2988,
"1101100100000011" when 2989,
"0001000010000111" when 2990,
"0011101100011101" when 2991,
"0011011101110001" when 2992,
"0000100001100011" when 2993,
"1101001011000110" when 2994,
"1100000010001011" when 2995,
"1101111111111000" when 2996,
"0001100001110101" when 2997,
"0011110111001111" when 2998,
"0011001011001100" when 2999,
"0000000000001001" when 3000,
"1100110101000000" when 3001,
"1100001000101100" when 3002,
"1110011101111010" when 3003,
"0001111111110111" when 3004,
"0011111101110010" when 3005,
"0010110101000111" when 3006,
"1111011110101111" when 3007,
"1100100010011000" when 3008,
"1100010011011100" when 3009,
"1110111101100111" when 3010,
"0010011011101110" when 3011,
"0011111111111111" when 3012,
"0010011011111101" when 3013,
"1110111101111001" when 3014,
"1100010011100011" when 3015,
"1100100010001111" when 3016,
"1111011110011101" when 3017,
"0010110100111010" when 3018,
"0011111101110101" when 3019,
"0010000000001000" when 3020,
"1110011110001011" when 3021,
"1100001000110001" when 3022,
"1100110100110100" when 3023,
"1111111111110111" when 3024,
"0011001011000000" when 3025,
"0011110111010100" when 3026,
"0001100010000110" when 3027,
"1110000000001001" when 3028,
"1100000010001110" when 3029,
"1101001010111001" when 3030,
"0000100001010001" when 3031,
"0011011101101000" when 3032,
"0011101100100100" when 3033,
"0001000010011001" when 3034,
"1101100100010010" when 3035,
"1100000000000001" when 3036,
"1101100100000011" when 3037,
"0001000010000111" when 3038,
"0011101100011101" when 3039,
"0011011101110001" when 3040,
"0000100001100011" when 3041,
"1101001011000110" when 3042,
"1100000010001011" when 3043,
"1101111111111000" when 3044,
"0001100001110101" when 3045,
"0011110111001111" when 3046,
"0011001011001100" when 3047,
"0000000000001001" when 3048,
"1100110101000000" when 3049,
"1100001000101100" when 3050,
"1110011101111010" when 3051,
"0001111111110111" when 3052,
"0011111101110010" when 3053,
"0010110101000111" when 3054,
"1111011110101111" when 3055,
"1100100010011000" when 3056,
"1100010011011100" when 3057,
"1110111101100111" when 3058,
"0010011011101110" when 3059,
"0011111111111111" when 3060,
"0010011011111101" when 3061,
"1110111101111001" when 3062,
"1100010011100011" when 3063,
"1100100010001111" when 3064,
"1111011110011100" when 3065,
"0010110100111010" when 3066,
"0011111101110101" when 3067,
"0010000000001000" when 3068,
"1110011110001011" when 3069,
"1100001000110001" when 3070,
"1100110100110100" when 3071,
"1111111111110111" when 3072,
"0011001011000000" when 3073,
"0011110111010100" when 3074,
"0001100010000110" when 3075,
"1110000000001001" when 3076,
"1100000010001110" when 3077,
"1101001010111000" when 3078,
"0000100001010001" when 3079,
"0011011101101000" when 3080,
"0011101100100100" when 3081,
"0001000010011001" when 3082,
"1101100100010010" when 3083,
"1100000000000001" when 3084,
"1101100100000011" when 3085,
"0001000010000111" when 3086,
"0011101100011101" when 3087,
"0011011101110001" when 3088,
"0000100001100100" when 3089,
"1101001011000110" when 3090,
"1100000010001011" when 3091,
"1101111111111000" when 3092,
"0001100001110100" when 3093,
"0011110111001111" when 3094,
"0011001011001100" when 3095,
"0000000000001001" when 3096,
"1100110101000000" when 3097,
"1100001000101100" when 3098,
"1110011101111010" when 3099,
"0001111111110111" when 3100,
"0011111101110010" when 3101,
"0010110101001000" when 3102,
"1111011110110000" when 3103,
"1100100010011000" when 3104,
"1100010011011100" when 3105,
"1110111101100111" when 3106,
"0010011011101110" when 3107,
"0011111111111111" when 3108,
"0010011011111101" when 3109,
"1110111101111001" when 3110,
"1100010011100011" when 3111,
"1100100010001111" when 3112,
"1111011110011100" when 3113,
"0010110100111010" when 3114,
"0011111101110101" when 3115,
"0010000000001000" when 3116,
"1110011110001100" when 3117,
"1100001000110001" when 3118,
"1100110100110100" when 3119,
"1111111111110111" when 3120,
"0011001011000000" when 3121,
"0011110111010100" when 3122,
"0001100010000110" when 3123,
"1110000000001001" when 3124,
"1100000010001110" when 3125,
"1101001010111000" when 3126,
"0000100001010000" when 3127,
"0011011101101000" when 3128,
"0011101100100100" when 3129,
"0001000010011001" when 3130,
"1101100100010010" when 3131,
"1100000000000001" when 3132,
"1101100100000011" when 3133,
"0001000010000111" when 3134,
"0011101100011101" when 3135,
"0011011101110001" when 3136,
"0000100001100100" when 3137,
"1101001011000110" when 3138,
"1100000010001011" when 3139,
"1101111111111000" when 3140,
"0001100001110100" when 3141,
"0011110111001111" when 3142,
"0011001011001100" when 3143,
"0000000000001001" when 3144,
"1100110101000000" when 3145,
"1100001000101100" when 3146,
"1110011101111010" when 3147,
"0001111111110111" when 3148,
"0011111101110010" when 3149,
"0010110101001000" when 3150,
"1111011110110000" when 3151,
"1100100010011000" when 3152,
"1100010011011100" when 3153,
"1110111101100110" when 3154,
"0010011011101110" when 3155,
"0011111111111111" when 3156,
"0010011011111101" when 3157,
"1110111101111010" when 3158,
"1100010011100011" when 3159,
"1100100010001111" when 3160,
"1111011110011100" when 3161,
"0010110100111010" when 3162,
"0011111101110101" when 3163,
"0010000000001000" when 3164,
"1110011110001100" when 3165,
"1100001000110001" when 3166,
"1100110100110100" when 3167,
"1111111111110111" when 3168,
"0011001011000000" when 3169,
"0011110111010100" when 3170,
"0001100010000111" when 3171,
"1110000000001001" when 3172,
"1100000010001110" when 3173,
"1101001010111000" when 3174,
"0000100001010000" when 3175,
"0011011101100111" when 3176,
"0011101100100100" when 3177,
"0001000010011010" when 3178,
"1101100100010010" when 3179,
"1100000000000001" when 3180,
"1101100100000011" when 3181,
"0001000010000110" when 3182,
"0011101100011101" when 3183,
"0011011101110001" when 3184,
"0000100001100100" when 3185,
"1101001011000110" when 3186,
"1100000010001011" when 3187,
"1101111111111000" when 3188,
"0001100001110100" when 3189,
"0011110111001111" when 3190,
"0011001011001100" when 3191,
"0000000000001001" when 3192,
"1100110101000000" when 3193,
"1100001000101100" when 3194,
"1110011101111001" when 3195,
"0001111111110111" when 3196,
"0011111101110010" when 3197,
"0010110101001000" when 3198,
"1111011110110000" when 3199,
"1100100010011001" when 3200,
"1100010011011100" when 3201,
"1110111101100110" when 3202,
"0010011011101110" when 3203,
"0011111111111111" when 3204,
"0010011011111101" when 3205,
"1110111101111010" when 3206,
"1100010011100011" when 3207,
"1100100010001111" when 3208,
"1111011110011100" when 3209,
"0010110100111010" when 3210,
"0011111101110101" when 3211,
"0010000000001000" when 3212,
"1110011110001100" when 3213,
"1100001000110001" when 3214,
"1100110100110100" when 3215,
"1111111111110110" when 3216,
"0011001011000000" when 3217,
"0011110111010100" when 3218,
"0001100010000111" when 3219,
"1110000000001001" when 3220,
"1100000010001110" when 3221,
"1101001010111000" when 3222,
"0000100001010000" when 3223,
"0011011101100111" when 3224,
"0011101100100100" when 3225,
"0001000010011010" when 3226,
"1101100100010011" when 3227,
"1100000000000001" when 3228,
"1101100100000011" when 3229,
"0001000010000110" when 3230,
"0011101100011100" when 3231,
"0011011101110010" when 3232,
"0000100001100100" when 3233,
"1101001011000110" when 3234,
"1100000010001011" when 3235,
"1101111111111000" when 3236,
"0001100001110100" when 3237,
"0011110111001111" when 3238,
"0011001011001100" when 3239,
"0000000000001010" when 3240,
"1100110101000000" when 3241,
"1100001000101100" when 3242,
"1110011101111001" when 3243,
"0001111111110111" when 3244,
"0011111101110010" when 3245,
"0010110101001000" when 3246,
"1111011110110000" when 3247,
"1100100010011001" when 3248,
"1100010011011100" when 3249,
"1110111101100110" when 3250,
"0010011011101101" when 3251,
"0011111111111111" when 3252,
"0010011011111110" when 3253,
"1110111101111010" when 3254,
"1100010011100100" when 3255,
"1100100010001110" when 3256,
"1111011110011100" when 3257,
"0010110100111010" when 3258,
"0011111101110101" when 3259,
"0010000000001000" when 3260,
"1110011110001100" when 3261,
"1100001000110001" when 3262,
"1100110100110100" when 3263,
"1111111111110110" when 3264,
"0011001011000000" when 3265,
"0011110111010100" when 3266,
"0001100010000111" when 3267,
"1110000000001001" when 3268,
"1100000010001110" when 3269,
"1101001010111000" when 3270,
"0000100001010000" when 3271,
"0011011101100111" when 3272,
"0011101100100100" when 3273,
"0001000010011010" when 3274,
"1101100100010011" when 3275,
"1100000000000001" when 3276,
"1101100100000010" when 3277,
"0001000010000110" when 3278,
"0011101100011100" when 3279,
"0011011101110010" when 3280,
"0000100001100100" when 3281,
"1101001011000111" when 3282,
"1100000010001011" when 3283,
"1101111111111000" when 3284,
"0001100001110100" when 3285,
"0011110111001111" when 3286,
"0011001011001100" when 3287,
"0000000000001010" when 3288,
"1100110101000000" when 3289,
"1100001000101100" when 3290,
"1110011101111001" when 3291,
"0001111111110111" when 3292,
"0011111101110010" when 3293,
"0010110101001000" when 3294,
"1111011110110000" when 3295,
"1100100010011001" when 3296,
"1100010011011100" when 3297,
"1110111101100110" when 3298,
"0010011011101101" when 3299,
"0011111111111111" when 3300,
"0010011011111110" when 3301,
"1110111101111010" when 3302,
"1100010011100100" when 3303,
"1100100010001110" when 3304,
"1111011110011100" when 3305,
"0010110100111001" when 3306,
"0011111101110101" when 3307,
"0010000000001000" when 3308,
"1110011110001100" when 3309,
"1100001000110001" when 3310,
"1100110100110100" when 3311,
"1111111111110110" when 3312,
"0011001010111111" when 3313,
"0011110111010100" when 3314,
"0001100010000111" when 3315,
"1110000000001001" when 3316,
"1100000010001110" when 3317,
"1101001010111000" when 3318,
"0000100001010000" when 3319,
"0011011101100111" when 3320,
"0011101100100100" when 3321,
"0001000010011010" when 3322,
"1101100100010011" when 3323,
"1100000000000001" when 3324,
"1101100100000010" when 3325,
"0001000010000110" when 3326,
"0011101100011100" when 3327,
"0011011101110010" when 3328,
"0000100001100100" when 3329,
"1101001011000111" when 3330,
"1100000010001011" when 3331,
"1101111111110111" when 3332,
"0001100001110100" when 3333,
"0011110111001111" when 3334,
"0011001011001100" when 3335,
"0000000000001010" when 3336,
"1100110101000001" when 3337,
"1100001000101100" when 3338,
"1110011101111001" when 3339,
"0001111111110110" when 3340,
"0011111101110010" when 3341,
"0010110101001000" when 3342,
"1111011110110000" when 3343,
"1100100010011001" when 3344,
"1100010011011100" when 3345,
"1110111101100110" when 3346,
"0010011011101101" when 3347,
"0011111111111111" when 3348,
"0010011011111110" when 3349,
"1110111101111010" when 3350,
"1100010011100100" when 3351,
"1100100010001110" when 3352,
"1111011110011100" when 3353,
"0010110100111001" when 3354,
"0011111101110101" when 3355,
"0010000000001001" when 3356,
"1110011110001100" when 3357,
"1100001000110001" when 3358,
"1100110100110100" when 3359,
"1111111111110110" when 3360,
"0011001010111111" when 3361,
"0011110111010100" when 3362,
"0001100010000111" when 3363,
"1110000000001010" when 3364,
"1100000010001110" when 3365,
"1101001010111000" when 3366,
"0000100001010000" when 3367,
"0011011101100111" when 3368,
"0011101100100100" when 3369,
"0001000010011010" when 3370,
"1101100100010011" when 3371,
"1100000000000001" when 3372,
"1101100100000010" when 3373,
"0001000010000110" when 3374,
"0011101100011100" when 3375,
"0011011101110010" when 3376,
"0000100001100100" when 3377,
"1101001011000111" when 3378,
"1100000010001011" when 3379,
"1101111111110111" when 3380,
"0001100001110100" when 3381,
"0011110111001110" when 3382,
"0011001011001100" when 3383,
"0000000000001010" when 3384,
"1100110101000001" when 3385,
"1100001000101100" when 3386,
"1110011101111001" when 3387,
"0001111111110110" when 3388,
"0011111101110010" when 3389,
"0010110101001000" when 3390,
"1111011110110000" when 3391,
"1100100010011001" when 3392,
"1100010011011100" when 3393,
"1110111101100110" when 3394,
"0010011011101101" when 3395,
"0011111111111111" when 3396,
"0010011011111110" when 3397,
"1110111101111010" when 3398,
"1100010011100100" when 3399,
"1100100010001110" when 3400,
"1111011110011011" when 3401,
"0010110100111001" when 3402,
"0011111101110101" when 3403,
"0010000000001001" when 3404,
"1110011110001100" when 3405,
"1100001000110010" when 3406,
"1100110100110100" when 3407,
"1111111111110110" when 3408,
"0011001010111111" when 3409,
"0011110111010100" when 3410,
"0001100010000111" when 3411,
"1110000000001010" when 3412,
"1100000010001110" when 3413,
"1101001010111000" when 3414,
"0000100001001111" when 3415,
"0011011101100111" when 3416,
"0011101100100100" when 3417,
"0001000010011010" when 3418,
"1101100100010011" when 3419,
"1100000000000001" when 3420,
"1101100100000010" when 3421,
"0001000010000110" when 3422,
"0011101100011100" when 3423,
"0011011101110010" when 3424,
"0000100001100101" when 3425,
"1101001011000111" when 3426,
"1100000010001011" when 3427,
"1101111111110111" when 3428,
"0001100001110011" when 3429,
"0011110111001110" when 3430,
"0011001011001100" when 3431,
"0000000000001010" when 3432,
"1100110101000001" when 3433,
"1100001000101100" when 3434,
"1110011101111001" when 3435,
"0001111111110110" when 3436,
"0011111101110010" when 3437,
"0010110101001000" when 3438,
"1111011110110001" when 3439,
"1100100010011001" when 3440,
"1100010011011100" when 3441,
"1110111101100110" when 3442,
"0010011011101101" when 3443,
"0011111111111111" when 3444,
"0010011011111110" when 3445,
"1110111101111010" when 3446,
"1100010011100100" when 3447,
"1100100010001110" when 3448,
"1111011110011011" when 3449,
"0010110100111001" when 3450,
"0011111101110101" when 3451,
"0010000000001001" when 3452,
"1110011110001101" when 3453,
"1100001000110010" when 3454,
"1100110100110100" when 3455,
"1111111111110110" when 3456,
"0011001010111111" when 3457,
"0011110111010100" when 3458,
"0001100010000111" when 3459,
"1110000000001010" when 3460,
"1100000010001110" when 3461,
"1101001010111000" when 3462,
"0000100001001111" when 3463,
"0011011101100111" when 3464,
"0011101100100100" when 3465,
"0001000010011010" when 3466,
"1101100100010011" when 3467,
"1100000000000001" when 3468,
"1101100100000010" when 3469,
"0001000010000110" when 3470,
"0011101100011100" when 3471,
"0011011101110010" when 3472,
"0000100001100101" when 3473,
"1101001011000111" when 3474,
"1100000010001011" when 3475,
"1101111111110111" when 3476,
"0001100001110011" when 3477,
"0011110111001110" when 3478,
"0011001011001100" when 3479,
"0000000000001010" when 3480,
"1100110101000001" when 3481,
"1100001000101100" when 3482,
"1110011101111001" when 3483,
"0001111111110110" when 3484,
"0011111101110010" when 3485,
"0010110101001000" when 3486,
"1111011110110001" when 3487,
"1100100010011001" when 3488,
"1100010011011011" when 3489,
"1110111101100101" when 3490,
"0010011011101101" when 3491,
"0011111111111111" when 3492,
"0010011011111110" when 3493,
"1110111101111011" when 3494,
"1100010011100100" when 3495,
"1100100010001110" when 3496,
"1111011110011011" when 3497,
"0010110100111001" when 3498,
"0011111101110101" when 3499,
"0010000000001001" when 3500,
"1110011110001101" when 3501,
"1100001000110010" when 3502,
"1100110100110100" when 3503,
"1111111111110110" when 3504,
"0011001010111111" when 3505,
"0011110111010100" when 3506,
"0001100010001000" when 3507,
"1110000000001010" when 3508,
"1100000010001110" when 3509,
"1101001010111000" when 3510,
"0000100001001111" when 3511,
"0011011101100111" when 3512,
"0011101100100101" when 3513,
"0001000010011011" when 3514,
"1101100100010011" when 3515,
"1100000000000001" when 3516,
"1101100100000010" when 3517,
"0001000010000101" when 3518,
"0011101100011100" when 3519,
"0011011101110010" when 3520,
"0000100001100101" when 3521,
"1101001011000111" when 3522,
"1100000010001011" when 3523,
"1101111111110111" when 3524,
"0001100001110011" when 3525,
"0011110111001110" when 3526,
"0011001011001101" when 3527,
"0000000000001011" when 3528,
"1100110101000001" when 3529,
"1100001000101100" when 3530,
"1110011101111000" when 3531,
"0001111111110110" when 3532,
"0011111101110010" when 3533,
"0010110101001001" when 3534,
"1111011110110001" when 3535,
"1100100010011001" when 3536,
"1100010011011011" when 3537,
"1110111101100101" when 3538,
"0010011011101101" when 3539,
"0011111111111111" when 3540,
"0010011011111110" when 3541,
"1110111101111011" when 3542,
"1100010011100100" when 3543,
"1100100010001110" when 3544,
"1111011110011011" when 3545,
"0010110100111001" when 3546,
"0011111101110101" when 3547,
"0010000000001001" when 3548,
"1110011110001101" when 3549,
"1100001000110010" when 3550,
"1100110100110011" when 3551,
"1111111111110101" when 3552,
"0011001010111111" when 3553,
"0011110111010100" when 3554,
"0001100010001000" when 3555,
"1110000000001010" when 3556,
"1100000010001110" when 3557,
"1101001010110111" when 3558,
"0000100001001111" when 3559,
"0011011101100111" when 3560,
"0011101100100101" when 3561,
"0001000010011011" when 3562,
"1101100100010011" when 3563,
"1100000000000001" when 3564,
"1101100100000010" when 3565,
"0001000010000101" when 3566,
"0011101100011100" when 3567,
"0011011101110010" when 3568,
"0000100001100101" when 3569,
"1101001011000111" when 3570,
"1100000010001011" when 3571,
"1101111111110111" when 3572,
"0001100001110011" when 3573,
"0011110111001110" when 3574,
"0011001011001101" when 3575,
"0000000000001011" when 3576,
"1100110101000001" when 3577,
"1100001000101100" when 3578,
"1110011101111000" when 3579,
"0001111111110110" when 3580,
"0011111101110010" when 3581,
"0010110101001001" when 3582,
"1111011110110001" when 3583,
"1100100010011001" when 3584,
"1100010011011011" when 3585,
"1110111101100101" when 3586,
"0010011011101101" when 3587,
"0011111111111111" when 3588,
"0010011011111110" when 3589,
"1110111101111011" when 3590,
"1100010011100100" when 3591,
"1100100010001110" when 3592,
"1111011110011011" when 3593,
"0010110100111001" when 3594,
"0011111101110101" when 3595,
"0010000000001001" when 3596,
"1110011110001101" when 3597,
"1100001000110010" when 3598,
"1100110100110011" when 3599,
"1111111111110101" when 3600,
"0011001010111111" when 3601,
"0011110111010100" when 3602,
"0001100010001000" when 3603,
"1110000000001010" when 3604,
"1100000010001110" when 3605,
"1101001010110111" when 3606,
"0000100001001111" when 3607,
"0011011101100111" when 3608,
"0011101100100101" when 3609,
"0001000010011011" when 3610,
"1101100100010100" when 3611,
"1100000000000001" when 3612,
"1101100100000010" when 3613,
"0001000010000101" when 3614,
"0011101100011100" when 3615,
"0011011101110010" when 3616,
"0000100001100101" when 3617,
"1101001011000111" when 3618,
"1100000010001011" when 3619,
"1101111111110111" when 3620,
"0001100001110011" when 3621,
"0011110111001110" when 3622,
"0011001011001101" when 3623,
"0000000000001011" when 3624,
"1100110101000001" when 3625,
"1100001000101100" when 3626,
"1110011101111000" when 3627,
"0001111111110110" when 3628,
"0011111101110010" when 3629,
"0010110101001001" when 3630,
"1111011110110001" when 3631,
"1100100010011001" when 3632,
"1100010011011011" when 3633,
"1110111101100101" when 3634,
"0010011011101100" when 3635,
"0011111111111111" when 3636,
"0010011011111110" when 3637,
"1110111101111011" when 3638,
"1100010011100100" when 3639,
"1100100010001110" when 3640,
"1111011110011011" when 3641,
"0010110100111001" when 3642,
"0011111101110101" when 3643,
"0010000000001001" when 3644,
"1110011110001101" when 3645,
"1100001000110010" when 3646,
"1100110100110011" when 3647,
"1111111111110101" when 3648,
"0011001010111111" when 3649,
"0011110111010100" when 3650,
"0001100010001000" when 3651,
"1110000000001010" when 3652,
"1100000010001110" when 3653,
"1101001010110111" when 3654,
"0000100001001111" when 3655,
"0011011101100111" when 3656,
"0011101100100101" when 3657,
"0001000010011011" when 3658,
"1101100100010100" when 3659,
"1100000000000001" when 3660,
"1101100100000001" when 3661,
"0001000010000101" when 3662,
"0011101100011100" when 3663,
"0011011101110010" when 3664,
"0000100001100101" when 3665,
"1101001011000111" when 3666,
"1100000010001011" when 3667,
"1101111111110111" when 3668,
"0001100001110011" when 3669,
"0011110111001110" when 3670,
"0011001011001101" when 3671,
"0000000000001011" when 3672,
"1100110101000001" when 3673,
"1100001000101100" when 3674,
"1110011101111000" when 3675,
"0001111111110110" when 3676,
"0011111101110010" when 3677,
"0010110101001001" when 3678,
"1111011110110001" when 3679,
"1100100010011001" when 3680,
"1100010011011011" when 3681,
"1110111101100101" when 3682,
"0010011011101100" when 3683,
"0011111111111111" when 3684,
"0010011011111111" when 3685,
"1110111101111011" when 3686,
"1100010011100100" when 3687,
"1100100010001110" when 3688,
"1111011110011011" when 3689,
"0010110100111001" when 3690,
"0011111101110101" when 3691,
"0010000000001001" when 3692,
"1110011110001101" when 3693,
"1100001000110010" when 3694,
"1100110100110011" when 3695,
"1111111111110101" when 3696,
"0011001010111111" when 3697,
"0011110111010100" when 3698,
"0001100010001000" when 3699,
"1110000000001011" when 3700,
"1100000010001110" when 3701,
"1101001010110111" when 3702,
"0000100001001111" when 3703,
"0011011101100111" when 3704,
"0011101100100101" when 3705,
"0001000010011011" when 3706,
"1101100100010100" when 3707,
"1100000000000001" when 3708,
"1101100100000001" when 3709,
"0001000010000101" when 3710,
"0011101100011100" when 3711,
"0011011101110010" when 3712,
"0000100001100110" when 3713,
"1101001011000111" when 3714,
"1100000010001011" when 3715,
"1101111111110110" when 3716,
"0001100001110011" when 3717,
"0011110111001110" when 3718,
"0011001011001101" when 3719,
"0000000000001011" when 3720,
"1100110101000001" when 3721,
"1100001000101100" when 3722,
"1110011101111000" when 3723,
"0001111111110101" when 3724,
"0011111101110010" when 3725,
"0010110101001001" when 3726,
"1111011110110010" when 3727,
"1100100010011001" when 3728,
"1100010011011011" when 3729,
"1110111101100101" when 3730,
"0010011011101100" when 3731,
"0011111111111111" when 3732,
"0010011011111111" when 3733,
"1110111101111011" when 3734,
"1100010011100100" when 3735,
"1100100010001110" when 3736,
"1111011110011010" when 3737,
"0010110100111000" when 3738,
"0011111101110101" when 3739,
"0010000000001010" when 3740,
"1110011110001101" when 3741,
"1100001000110010" when 3742,
"1100110100110011" when 3743,
"1111111111110101" when 3744,
"0011001010111111" when 3745,
"0011110111010100" when 3746,
"0001100010001000" when 3747,
"1110000000001011" when 3748,
"1100000010001110" when 3749,
"1101001010110111" when 3750,
"0000100001001110" when 3751,
"0011011101100111" when 3752,
"0011101100100101" when 3753,
"0001000010011011" when 3754,
"1101100100010100" when 3755,
"1100000000000001" when 3756,
"1101100100000001" when 3757,
"0001000010000101" when 3758,
"0011101100011100" when 3759,
"0011011101110010" when 3760,
"0000100001100110" when 3761,
"1101001011001000" when 3762,
"1100000010001011" when 3763,
"1101111111110110" when 3764,
"0001100001110011" when 3765,
"0011110111001110" when 3766,
"0011001011001101" when 3767,
"0000000000001011" when 3768,
"1100110101000001" when 3769,
"1100001000101100" when 3770,
"1110011101111000" when 3771,
"0001111111110101" when 3772,
"0011111101110010" when 3773,
"0010110101001001" when 3774,
"1111011110110010" when 3775,
"1100100010011001" when 3776,
"1100010011011011" when 3777,
"1110111101100101" when 3778,
"0010011011101100" when 3779,
"0011111111111111" when 3780,
"0010011011111111" when 3781,
"1110111101111011" when 3782,
"1100010011100100" when 3783,
"1100100010001110" when 3784,
"1111011110011010" when 3785,
"0010110100111000" when 3786,
"0011111101110101" when 3787,
"0010000000001010" when 3788,
"1110011110001110" when 3789,
"1100001000110010" when 3790,
"1100110100110011" when 3791,
"1111111111110101" when 3792,
"0011001010111111" when 3793,
"0011110111010100" when 3794,
"0001100010001000" when 3795,
"1110000000001011" when 3796,
"1100000010001110" when 3797,
"1101001010110111" when 3798,
"0000100001001110" when 3799,
"0011011101100111" when 3800,
"0011101100100101" when 3801,
"0001000010011011" when 3802,
"1101100100010100" when 3803,
"1100000000000001" when 3804,
"1101100100000001" when 3805,
"0001000010000101" when 3806,
"0011101100011100" when 3807,
"0011011101110010" when 3808,
"0000100001100110" when 3809,
"1101001011001000" when 3810,
"1100000010001011" when 3811,
"1101111111110110" when 3812,
"0001100001110010" when 3813,
"0011110111001110" when 3814,
"0011001011001101" when 3815,
"0000000000001011" when 3816,
"1100110101000001" when 3817,
"1100001000101100" when 3818,
"1110011101111000" when 3819,
"0001111111110101" when 3820,
"0011111101110010" when 3821,
"0010110101001001" when 3822,
"1111011110110010" when 3823,
"1100100010011010" when 3824,
"1100010011011011" when 3825,
"1110111101100100" when 3826,
"0010011011101100" when 3827,
"0011111111111111" when 3828,
"0010011011111111" when 3829,
"1110111101111100" when 3830,
"1100010011100100" when 3831,
"1100100010001110" when 3832,
"1111011110011010" when 3833,
"0010110100111000" when 3834,
"0011111101110101" when 3835,
"0010000000001010" when 3836,
"1110011110001110" when 3837,
"1100001000110010" when 3838,
"1100110100110011" when 3839,
"1111111111110101" when 3840,
"0011001010111110" when 3841,
"0011110111010100" when 3842,
"0001100010001000" when 3843,
"1110000000001011" when 3844,
"1100000010001110" when 3845,
"1101001010110111" when 3846,
"0000100001001110" when 3847,
"0011011101100110" when 3848,
"0011101100100101" when 3849,
"0001000010011100" when 3850,
"1101100100010100" when 3851,
"1100000000000001" when 3852,
"1101100100000001" when 3853,
"0001000010000100" when 3854,
"0011101100011100" when 3855,
"0011011101110010" when 3856,
"0000100001100110" when 3857,
"1101001011001000" when 3858,
"1100000010001011" when 3859,
"1101111111110110" when 3860,
"0001100001110010" when 3861,
"0011110111001110" when 3862,
"0011001011001101" when 3863,
"0000000000001100" when 3864,
"1100110101000010" when 3865,
"1100001000101100" when 3866,
"1110011101110111" when 3867,
"0001111111110101" when 3868,
"0011111101110010" when 3869,
"0010110101001001" when 3870,
"1111011110110010" when 3871,
"1100100010011010" when 3872,
"1100010011011011" when 3873,
"1110111101100100" when 3874,
"0010011011101100" when 3875,
"0011111111111111" when 3876,
"0010011011111111" when 3877,
"1110111101111100" when 3878,
"1100010011100100" when 3879,
"1100100010001101" when 3880,
"1111011110011010" when 3881,
"0010110100111000" when 3882,
"0011111101110101" when 3883,
"0010000000001010" when 3884,
"1110011110001110" when 3885,
"1100001000110010" when 3886,
"1100110100110011" when 3887,
"1111111111110100" when 3888,
"0011001010111110" when 3889,
"0011110111010100" when 3890,
"0001100010001001" when 3891,
"1110000000001011" when 3892,
"1100000010001110" when 3893,
"1101001010110111" when 3894,
"0000100001001110" when 3895,
"0011011101100110" when 3896,
"0011101100100101" when 3897,
"0001000010011100" when 3898,
"1101100100010100" when 3899,
"1100000000000001" when 3900,
"1101100100000001" when 3901,
"0001000010000100" when 3902,
"0011101100011100" when 3903,
"0011011101110011" when 3904,
"0000100001100110" when 3905,
"1101001011001000" when 3906,
"1100000010001011" when 3907,
"1101111111110110" when 3908,
"0001100001110010" when 3909,
"0011110111001110" when 3910,
"0011001011001101" when 3911,
"0000000000001100" when 3912,
"1100110101000010" when 3913,
"1100001000101100" when 3914,
"1110011101110111" when 3915,
"0001111111110101" when 3916,
"0011111101110010" when 3917,
"0010110101001001" when 3918,
"1111011110110010" when 3919,
"1100100010011010" when 3920,
"1100010011011011" when 3921,
"1110111101100100" when 3922,
"0010011011101100" when 3923,
"0011111111111111" when 3924,
"0010011011111111" when 3925,
"1110111101111100" when 3926,
"1100010011100100" when 3927,
"1100100010001101" when 3928,
"1111011110011010" when 3929,
"0010110100111000" when 3930,
"0011111101110101" when 3931,
"0010000000001010" when 3932,
"1110011110001110" when 3933,
"1100001000110010" when 3934,
"1100110100110011" when 3935,
"1111111111110100" when 3936,
"0011001010111110" when 3937,
"0011110111010100" when 3938,
"0001100010001001" when 3939,
"1110000000001011" when 3940,
"1100000010001110" when 3941,
"1101001010110111" when 3942,
"0000100001001110" when 3943,
"0011011101100110" when 3944,
"0011101100100101" when 3945,
"0001000010011100" when 3946,
"1101100100010100" when 3947,
"1100000000000001" when 3948,
"1101100100000001" when 3949,
"0001000010000100" when 3950,
"0011101100011100" when 3951,
"0011011101110011" when 3952,
"0000100001100110" when 3953,
"1101001011001000" when 3954,
"1100000010001011" when 3955,
"1101111111110110" when 3956,
"0001100001110010" when 3957,
"0011110111001110" when 3958,
"0011001011001101" when 3959,
"0000000000001100" when 3960,
"1100110101000010" when 3961,
"1100001000101100" when 3962,
"1110011101110111" when 3963,
"0001111111110101" when 3964,
"0011111101110010" when 3965,
"0010110101001001" when 3966,
"1111011110110010" when 3967,
"1100100010011010" when 3968,
"1100010011011011" when 3969,
"1110111101100100" when 3970,
"0010011011101100" when 3971,
"0011111111111111" when 3972,
"0010011011111111" when 3973,
"1110111101111100" when 3974,
"1100010011100100" when 3975,
"1100100010001101" when 3976,
"1111011110011010" when 3977,
"0010110100111000" when 3978,
"0011111101110101" when 3979,
"0010000000001010" when 3980,
"1110011110001110" when 3981,
"1100001000110010" when 3982,
"1100110100110011" when 3983,
"1111111111110100" when 3984,
"0011001010111110" when 3985,
"0011110111010100" when 3986,
"0001100010001001" when 3987,
"1110000000001011" when 3988,
"1100000010001110" when 3989,
"1101001010110110" when 3990,
"0000100001001110" when 3991,
"0011011101100110" when 3992,
"0011101100100101" when 3993,
"0001000010011100" when 3994,
"1101100100010100" when 3995,
"1100000000000001" when 3996,
"1101100100000001" when 3997,
"0001000010000100" when 3998,
"0011101100011100" when 3999,
"0011011101110011" when 4000,
"0000100001100110" when 4001,
"1101001011001000" when 4002,
"1100000010001011" when 4003,
"1101111111110110" when 4004,
"0001100001110010" when 4005,
"0011110111001110" when 4006,
"0011001011001101" when 4007,
"0000000000001100" when 4008,
"1100110101000010" when 4009,
"1100001000101100" when 4010,
"1110011101110111" when 4011,
"0001111111110101" when 4012,
"0011111101110010" when 4013,
"0010110101001010" when 4014,
"1111011110110010" when 4015,
"1100100010011010" when 4016,
"1100010011011011" when 4017,
"1110111101100100" when 4018,
"0010011011101011" when 4019,
"0011111111111111" when 4020,
"0010011011111111" when 4021,
"1110111101111100" when 4022,
"1100010011100100" when 4023,
"1100100010001101" when 4024,
"1111011110011001" when 4025,
"0010110100111000" when 4026,
"0011111101110101" when 4027,
"0010000000001010" when 4028,
"1110011110001110" when 4029,
"1100001000110010" when 4030,
"1100110100110011" when 4031,
"1111111111110100" when 4032,
"0011001010111110" when 4033,
"0011110111010100" when 4034,
"0001100010001001" when 4035,
"1110000000001011" when 4036,
"1100000010001110" when 4037,
"1101001010110110" when 4038,
"0000100001001110" when 4039,
"0011011101100110" when 4040,
"0011101100100101" when 4041,
"0001000010011100" when 4042,
"1101100100010101" when 4043,
"1100000000000001" when 4044,
"1101100100000001" when 4045,
"0001000010000100" when 4046,
"0011101100011100" when 4047,
"0011011101110011" when 4048,
"0000100001100111" when 4049,
"1101001011001000" when 4050,
"1100000010001011" when 4051,
"1101111111110110" when 4052,
"0001100001110010" when 4053,
"0011110111001110" when 4054,
"0011001011001110" when 4055,
"0000000000001100" when 4056,
"1100110101000010" when 4057,
"1100001000101011" when 4058,
"1110011101110111" when 4059,
"0001111111110101" when 4060,
"0011111101110010" when 4061,
"0010110101001010" when 4062,
"1111011110110011" when 4063,
"1100100010011010" when 4064,
"1100010011011011" when 4065,
"1110111101100100" when 4066,
"0010011011101011" when 4067,
"0011111111111111" when 4068,
"0010011100000000" when 4069,
"1110111101111100" when 4070,
"1100010011100101" when 4071,
"1100100010001101" when 4072,
"1111011110011001" when 4073,
"0010110100111000" when 4074,
"0011111101110101" when 4075,
"0010000000001011" when 4076,
"1110011110001110" when 4077,
"1100001000110010" when 4078,
"1100110100110010" when 4079,
"1111111111110100" when 4080,
"0011001010111110" when 4081,
"0011110111010101" when 4082,
"0001100010001001" when 4083,
"1110000000001100" when 4084,
"1100000010001110" when 4085,
"1101001010110110" when 4086,
"0000100001001101" when 4087,
"0011011101100110" when 4088,
"0011101100100101" when 4089,
"0001000010011100" when 4090,
"1101100100010101" when 4091,
"1100000000000001" when 4092,
"1101100100000000" when 4093,
"0001000010000100" when 4094,
"0011101100011011" when 4095,
"0011011101110011" when 4096,
"0000100001100111" when 4097,
"1101001011001000" when 4098,
"1100000010001011" when 4099,
"1101111111110101" when 4100,
"0001100001110010" when 4101,
"0011110111001110" when 4102,
"0011001011001110" when 4103,
"0000000000001100" when 4104,
"1100110101000010" when 4105,
"1100001000101011" when 4106,
"1110011101110111" when 4107,
"0001111111110100" when 4108,
"0011111101110010" when 4109,
"0010110101001010" when 4110,
"1111011110110011" when 4111,
"1100100010011010" when 4112,
"1100010011011011" when 4113,
"1110111101100100" when 4114,
"0010011011101011" when 4115,
"0011111111111111" when 4116,
"0010011100000000" when 4117,
"1110111101111100" when 4118,
"1100010011100101" when 4119,
"1100100010001101" when 4120,
"1111011110011001" when 4121,
"0010110100111000" when 4122,
"0011111101110101" when 4123,
"0010000000001011" when 4124,
"1110011110001111" when 4125,
"1100001000110010" when 4126,
"1100110100110010" when 4127,
"1111111111110100" when 4128,
"0011001010111110" when 4129,
"0011110111010101" when 4130,
"0001100010001001" when 4131,
"1110000000001100" when 4132,
"1100000010001110" when 4133,
"1101001010110110" when 4134,
"0000100001001101" when 4135,
"0011011101100110" when 4136,
"0011101100100101" when 4137,
"0001000010011100" when 4138,
"1101100100010101" when 4139,
"1100000000000001" when 4140,
"1101100100000000" when 4141,
"0001000010000011" when 4142,
"0011101100011011" when 4143,
"0011011101110011" when 4144,
"0000100001100111" when 4145,
"1101001011001000" when 4146,
"1100000010001011" when 4147,
"1101111111110101" when 4148,
"0001100001110001" when 4149,
"0011110111001110" when 4150,
"0011001011001110" when 4151,
"0000000000001100" when 4152,
"1100110101000010" when 4153,
"1100001000101011" when 4154,
"1110011101110111" when 4155,
"0001111111110100" when 4156,
"0011111101110010" when 4157,
"0010110101001010" when 4158,
"1111011110110011" when 4159,
"1100100010011010" when 4160,
"1100010011011011" when 4161,
"1110111101100011" when 4162,
"0010011011101011" when 4163,
"0011111111111111" when 4164,
"0010011100000000" when 4165,
"1110111101111101" when 4166,
"1100010011100101" when 4167,
"1100100010001101" when 4168,
"1111011110011001" when 4169,
"0010110100111000" when 4170,
"0011111101110101" when 4171,
"0010000000001011" when 4172,
"1110011110001111" when 4173,
"1100001000110010" when 4174,
"1100110100110010" when 4175,
"1111111111110011" when 4176,
"0011001010111110" when 4177,
"0011110111010101" when 4178,
"0001100010001001" when 4179,
"1110000000001100" when 4180,
"1100000010001110" when 4181,
"1101001010110110" when 4182,
"0000100001001101" when 4183,
"0011011101100110" when 4184,
"0011101100100101" when 4185,
"0001000010011101" when 4186,
"1101100100010101" when 4187,
"1100000000000001" when 4188,
"1101100100000000" when 4189,
"0001000010000011" when 4190,
"0011101100011011" when 4191,
"0011011101110011" when 4192,
"0000100001100111" when 4193,
"1101001011001001" when 4194,
"1100000010001011" when 4195,
"1101111111110101" when 4196,
"0001100001110001" when 4197,
"0011110111001110" when 4198,
"0011001011001110" when 4199,
"0000000000001101" when 4200,
"1100110101000010" when 4201,
"1100001000101011" when 4202,
"1110011101110110" when 4203,
"0001111111110100" when 4204,
"0011111101110010" when 4205,
"0010110101001010" when 4206,
"1111011110110011" when 4207,
"1100100010011010" when 4208,
"1100010011011011" when 4209,
"1110111101100011" when 4210,
"0010011011101011" when 4211,
"0011111111111111" when 4212,
"0010011100000000" when 4213,
"1110111101111101" when 4214,
"1100010011100101" when 4215,
"1100100010001101" when 4216,
"1111011110011001" when 4217,
"0010110100110111" when 4218,
"0011111101110101" when 4219,
"0010000000001011" when 4220,
"1110011110001111" when 4221,
"1100001000110010" when 4222,
"1100110100110010" when 4223,
"1111111111110011" when 4224,
"0011001010111110" when 4225,
"0011110111010101" when 4226,
"0001100010001010" when 4227,
"1110000000001100" when 4228,
"1100000010001110" when 4229,
"1101001010110110" when 4230,
"0000100001001101" when 4231,
"0011011101100110" when 4232,
"0011101100100101" when 4233,
"0001000010011101" when 4234,
"1101100100010101" when 4235,
"1100000000000001" when 4236,
"1101100100000000" when 4237,
"0001000010000011" when 4238,
"0011101100011011" when 4239,
"0011011101110011" when 4240,
"0000100001100111" when 4241,
"1101001011001001" when 4242,
"1100000010001011" when 4243,
"1101111111110101" when 4244,
"0001100001110001" when 4245,
"0011110111001110" when 4246,
"0011001011001110" when 4247,
"0000000000001101" when 4248,
"1100110101000010" when 4249,
"1100001000101011" when 4250,
"1110011101110110" when 4251,
"0001111111110100" when 4252,
"0011111101110010" when 4253,
"0010110101001010" when 4254,
"1111011110110011" when 4255,
"1100100010011010" when 4256,
"1100010011011011" when 4257,
"1110111101100011" when 4258,
"0010011011101011" when 4259,
"0011111111111111" when 4260,
"0010011100000000" when 4261,
"1110111101111101" when 4262,
"1100010011100101" when 4263,
"1100100010001101" when 4264,
"1111011110011001" when 4265,
"0010110100110111" when 4266,
"0011111101110101" when 4267,
"0010000000001011" when 4268,
"1110011110001111" when 4269,
"1100001000110010" when 4270,
"1100110100110010" when 4271,
"1111111111110011" when 4272,
"0011001010111110" when 4273,
"0011110111010101" when 4274,
"0001100010001010" when 4275,
"1110000000001100" when 4276,
"1100000010001110" when 4277,
"1101001010110110" when 4278,
"0000100001001101" when 4279,
"0011011101100110" when 4280,
"0011101100100101" when 4281,
"0001000010011101" when 4282,
"1101100100010101" when 4283,
"1100000000000001" when 4284,
"1101100100000000" when 4285,
"0001000010000011" when 4286,
"0011101100011011" when 4287,
"0011011101110011" when 4288,
"0000100001100111" when 4289,
"1101001011001001" when 4290,
"1100000010001011" when 4291,
"1101111111110101" when 4292,
"0001100001110001" when 4293,
"0011110111001110" when 4294,
"0011001011001110" when 4295,
"0000000000001101" when 4296,
"1100110101000010" when 4297,
"1100001000101011" when 4298,
"1110011101110110" when 4299,
"0001111111110100" when 4300,
"0011111101110010" when 4301,
"0010110101001010" when 4302,
"1111011110110011" when 4303,
"1100100010011010" when 4304,
"1100010011011011" when 4305,
"1110111101100011" when 4306,
"0010011011101011" when 4307,
"0011111111111111" when 4308,
"0010011100000000" when 4309,
"1110111101111101" when 4310,
"1100010011100101" when 4311,
"1100100010001101" when 4312,
"1111011110011001" when 4313,
"0010110100110111" when 4314,
"0011111101110101" when 4315,
"0010000000001011" when 4316,
"1110011110001111" when 4317,
"1100001000110010" when 4318,
"1100110100110010" when 4319,
"1111111111110011" when 4320,
"0011001010111110" when 4321,
"0011110111010101" when 4322,
"0001100010001010" when 4323,
"1110000000001100" when 4324,
"1100000010001110" when 4325,
"1101001010110110" when 4326,
"0000100001001101" when 4327,
"0011011101100110" when 4328,
"0011101100100110" when 4329,
"0001000010011101" when 4330,
"1101100100010101" when 4331,
"1100000000000001" when 4332,
"1101100100000000" when 4333,
"0001000010000011" when 4334,
"0011101100011011" when 4335,
"0011011101110011" when 4336,
"0000100001100111" when 4337,
"1101001011001001" when 4338,
"1100000010001011" when 4339,
"1101111111110101" when 4340,
"0001100001110001" when 4341,
"0011110111001110" when 4342,
"0011001011001110" when 4343,
"0000000000001101" when 4344,
"1100110101000010" when 4345,
"1100001000101011" when 4346,
"1110011101110110" when 4347,
"0001111111110100" when 4348,
"0011111101110010" when 4349,
"0010110101001010" when 4350,
"1111011110110011" when 4351,
"1100100010011010" when 4352,
"1100010011011010" when 4353,
"1110111101100011" when 4354,
"0010011011101011" when 4355,
"0011111111111111" when 4356,
"0010011100000000" when 4357,
"1110111101111101" when 4358,
"1100010011100101" when 4359,
"1100100010001101" when 4360,
"1111011110011000" when 4361,
"0010110100110111" when 4362,
"0011111101110101" when 4363,
"0010000000001011" when 4364,
"1110011110001111" when 4365,
"1100001000110010" when 4366,
"1100110100110010" when 4367,
"1111111111110011" when 4368,
"0011001010111101" when 4369,
"0011110111010101" when 4370,
"0001100010001010" when 4371,
"1110000000001100" when 4372,
"1100000010001110" when 4373,
"1101001010110110" when 4374,
"0000100001001100" when 4375,
"0011011101100110" when 4376,
"0011101100100110" when 4377,
"0001000010011101" when 4378,
"1101100100010101" when 4379,
"1100000000000001" when 4380,
"1101100100000000" when 4381,
"0001000010000011" when 4382,
"0011101100011011" when 4383,
"0011011101110011" when 4384,
"0000100001101000" when 4385,
"1101001011001001" when 4386,
"1100000010001011" when 4387,
"1101111111110101" when 4388,
"0001100001110001" when 4389,
"0011110111001110" when 4390,
"0011001011001110" when 4391,
"0000000000001101" when 4392,
"1100110101000011" when 4393,
"1100001000101011" when 4394,
"1110011101110110" when 4395,
"0001111111110100" when 4396,
"0011111101110010" when 4397,
"0010110101001010" when 4398,
"1111011110110100" when 4399,
"1100100010011010" when 4400,
"1100010011011010" when 4401,
"1110111101100011" when 4402,
"0010011011101011" when 4403,
"0011111111111111" when 4404,
"0010011100000000" when 4405,
"1110111101111101" when 4406,
"1100010011100101" when 4407,
"1100100010001101" when 4408,
"1111011110011000" when 4409,
"0010110100110111" when 4410,
"0011111101110101" when 4411,
"0010000000001011" when 4412,
"1110011110001111" when 4413,
"1100001000110010" when 4414,
"1100110100110010" when 4415,
"1111111111110011" when 4416,
"0011001010111101" when 4417,
"0011110111010101" when 4418,
"0001100010001010" when 4419,
"1110000000001100" when 4420,
"1100000010001110" when 4421,
"1101001010110110" when 4422,
"0000100001001100" when 4423,
"0011011101100110" when 4424,
"0011101100100110" when 4425,
"0001000010011101" when 4426,
"1101100100010110" when 4427,
"1100000000000001" when 4428,
"1101100100000000" when 4429,
"0001000010000011" when 4430,
"0011101100011011" when 4431,
"0011011101110011" when 4432,
"0000100001101000" when 4433,
"1101001011001001" when 4434,
"1100000010001011" when 4435,
"1101111111110101" when 4436,
"0001100001110001" when 4437,
"0011110111001110" when 4438,
"0011001011001110" when 4439,
"0000000000001101" when 4440,
"1100110101000011" when 4441,
"1100001000101011" when 4442,
"1110011101110110" when 4443,
"0001111111110011" when 4444,
"0011111101110010" when 4445,
"0010110101001011" when 4446,
"1111011110110100" when 4447,
"1100100010011010" when 4448,
"1100010011011010" when 4449,
"1110111101100011" when 4450,
"0010011011101010" when 4451,
"0011111111111111" when 4452,
"0010011100000000" when 4453,
"1110111101111101" when 4454,
"1100010011100101" when 4455,
"1100100010001101" when 4456,
"1111011110011000" when 4457,
"0010110100110111" when 4458,
"0011111101110101" when 4459,
"0010000000001100" when 4460,
"1110011110001111" when 4461,
"1100001000110010" when 4462,
"1100110100110010" when 4463,
"1111111111110011" when 4464,
"0011001010111101" when 4465,
"0011110111010101" when 4466,
"0001100010001010" when 4467,
"1110000000001101" when 4468,
"1100000010001110" when 4469,
"1101001010110101" when 4470,
"0000100001001100" when 4471,
"0011011101100101" when 4472,
"0011101100100110" when 4473,
"0001000010011101" when 4474,
"1101100100010110" when 4475,
"1100000000000001" when 4476,
"1101100011111111" when 4477,
"0001000010000010" when 4478,
"0011101100011011" when 4479,
"0011011101110011" when 4480,
"0000100001101000" when 4481,
"1101001011001001" when 4482,
"1100000010001011" when 4483,
"1101111111110100" when 4484,
"0001100001110000" when 4485,
"0011110111001110" when 4486,
"0011001011001110" when 4487,
"0000000000001110" when 4488,
"1100110101000011" when 4489,
"1100001000101011" when 4490,
"1110011101110110" when 4491,
"0001111111110011" when 4492,
"0011111101110001" when 4493,
"0010110101001011" when 4494,
"1111011110110100" when 4495,
"1100100010011011" when 4496,
"1100010011011010" when 4497,
"1110111101100010" when 4498,
"0010011011101010" when 4499,
"0011111111111111" when 4500,
"0010011100000001" when 4501,
"1110111101111110" when 4502,
"1100010011100101" when 4503,
"1100100010001101" when 4504,
"1111011110011000" when 4505,
"0010110100110111" when 4506,
"0011111101110101" when 4507,
"0010000000001100" when 4508,
"1110011110010000" when 4509,
"1100001000110010" when 4510,
"1100110100110010" when 4511,
"1111111111110010" when 4512,
"0011001010111101" when 4513,
"0011110111010101" when 4514,
"0001100010001010" when 4515,
"1110000000001101" when 4516,
"1100000010001111" when 4517,
"1101001010110101" when 4518,
"0000100001001100" when 4519,
"0011011101100101" when 4520,
"0011101100100110" when 4521,
"0001000010011110" when 4522,
"1101100100010110" when 4523,
"1100000000000001" when 4524,
"1101100011111111" when 4525,
"0001000010000010" when 4526,
"0011101100011011" when 4527,
"0011011101110100" when 4528,
"0000100001101000" when 4529,
"1101001011001001" when 4530,
"1100000010001011" when 4531,
"1101111111110100" when 4532,
"0001100001110000" when 4533,
"0011110111001110" when 4534,
"0011001011001110" when 4535,
"0000000000001110" when 4536,
"1100110101000011" when 4537,
"1100001000101011" when 4538,
"1110011101110110" when 4539,
"0001111111110011" when 4540,
"0011111101110001" when 4541,
"0010110101001011" when 4542,
"1111011110110100" when 4543,
"1100100010011011" when 4544,
"1100010011011010" when 4545,
"1110111101100010" when 4546,
"0010011011101010" when 4547,
"0011111111111111" when 4548,
"0010011100000001" when 4549,
"1110111101111110" when 4550,
"1100010011100101" when 4551,
"1100100010001100" when 4552,
"1111011110011000" when 4553,
"0010110100110111" when 4554,
"0011111101110101" when 4555,
"0010000000001100" when 4556,
"1110011110010000" when 4557,
"1100001000110010" when 4558,
"1100110100110010" when 4559,
"1111111111110010" when 4560,
"0011001010111101" when 4561,
"0011110111010101" when 4562,
"0001100010001011" when 4563,
"1110000000001101" when 4564,
"1100000010001111" when 4565,
"1101001010110101" when 4566,
"0000100001001100" when 4567,
"0011011101100101" when 4568,
"0011101100100110" when 4569,
"0001000010011110" when 4570,
"1101100100010110" when 4571,
"1100000000000001" when 4572,
"1101100011111111" when 4573,
"0001000010000010" when 4574,
"0011101100011011" when 4575,
"0011011101110100" when 4576,
"0000100001101000" when 4577,
"1101001011001001" when 4578,
"1100000010001011" when 4579,
"1101111111110100" when 4580,
"0001100001110000" when 4581,
"0011110111001110" when 4582,
"0011001011001111" when 4583,
"0000000000001110" when 4584,
"1100110101000011" when 4585,
"1100001000101011" when 4586,
"1110011101110101" when 4587,
"0001111111110011" when 4588,
"0011111101110001" when 4589,
"0010110101001011" when 4590,
"1111011110110100" when 4591,
"1100100010011011" when 4592,
"1100010011011010" when 4593,
"1110111101100010" when 4594,
"0010011011101010" when 4595,
"0011111111111111" when 4596,
"0010011100000001" when 4597,
"1110111101111110" when 4598,
"1100010011100101" when 4599,
"1100100010001100" when 4600,
"1111011110011000" when 4601,
"0010110100110111" when 4602,
"0011111101110101" when 4603,
"0010000000001100" when 4604,
"1110011110010000" when 4605,
"1100001000110011" when 4606,
"1100110100110001" when 4607,
"1111111111110010" when 4608,
"0011001010111101" when 4609,
"0011110111010101" when 4610,
"0001100010001011" when 4611,
"1110000000001101" when 4612,
"1100000010001111" when 4613,
"1101001010110101" when 4614,
"0000100001001100" when 4615,
"0011011101100101" when 4616,
"0011101100100110" when 4617,
"0001000010011110" when 4618,
"1101100100010110" when 4619,
"1100000000000001" when 4620,
"1101100011111111" when 4621,
"0001000010000010" when 4622,
"0011101100011011" when 4623,
"0011011101110100" when 4624,
"0000100001101000" when 4625,
"1101001011001001" when 4626,
"1100000010001011" when 4627,
"1101111111110100" when 4628,
"0001100001110000" when 4629,
"0011110111001101" when 4630,
"0011001011001111" when 4631,
"0000000000001110" when 4632,
"1100110101000011" when 4633,
"1100001000101011" when 4634,
"1110011101110101" when 4635,
"0001111111110011" when 4636,
"0011111101110001" when 4637,
"0010110101001011" when 4638,
"1111011110110100" when 4639,
"1100100010011011" when 4640,
"1100010011011010" when 4641,
"1110111101100010" when 4642,
"0010011011101010" when 4643,
"0011111111111111" when 4644,
"0010011100000001" when 4645,
"1110111101111110" when 4646,
"1100010011100101" when 4647,
"1100100010001100" when 4648,
"1111011110011000" when 4649,
"0010110100110110" when 4650,
"0011111101110101" when 4651,
"0010000000001100" when 4652,
"1110011110010000" when 4653,
"1100001000110011" when 4654,
"1100110100110001" when 4655,
"1111111111110010" when 4656,
"0011001010111101" when 4657,
"0011110111010101" when 4658,
"0001100010001011" when 4659,
"1110000000001101" when 4660,
"1100000010001111" when 4661,
"1101001010110101" when 4662,
"0000100001001100" when 4663,
"0011011101100101" when 4664,
"0011101100100110" when 4665,
"0001000010011110" when 4666,
"1101100100010110" when 4667,
"1100000000000001" when 4668,
"1101100011111111" when 4669,
"0001000010000010" when 4670,
"0011101100011011" when 4671,
"0011011101110100" when 4672,
"0000100001101001" when 4673,
"1101001011001010" when 4674,
"1100000010001011" when 4675,
"1101111111110100" when 4676,
"0001100001110000" when 4677,
"0011110111001101" when 4678,
"0011001011001111" when 4679,
"0000000000001110" when 4680,
"1100110101000011" when 4681,
"1100001000101011" when 4682,
"1110011101110101" when 4683,
"0001111111110011" when 4684,
"0011111101110001" when 4685,
"0010110101001011" when 4686,
"1111011110110100" when 4687,
"1100100010011011" when 4688,
"1100010011011010" when 4689,
"1110111101100010" when 4690,
"0010011011101010" when 4691,
"0011111111111111" when 4692,
"0010011100000001" when 4693,
"1110111101111110" when 4694,
"1100010011100101" when 4695,
"1100100010001100" when 4696,
"1111011110010111" when 4697,
"0010110100110110" when 4698,
"0011111101110101" when 4699,
"0010000000001100" when 4700,
"1110011110010000" when 4701,
"1100001000110011" when 4702,
"1100110100110001" when 4703,
"1111111111110010" when 4704,
"0011001010111101" when 4705,
"0011110111010101" when 4706,
"0001100010001011" when 4707,
"1110000000001101" when 4708,
"1100000010001111" when 4709,
"1101001010110101" when 4710,
"0000100001001011" when 4711,
"0011011101100101" when 4712,
"0011101100100110" when 4713,
"0001000010011110" when 4714,
"1101100100010110" when 4715,
"1100000000000001" when 4716,
"1101100011111111" when 4717,
"0001000010000010" when 4718,
"0011101100011011" when 4719,
"0011011101110100" when 4720,
"0000100001101001" when 4721,
"1101001011001010" when 4722,
"1100000010001011" when 4723,
"1101111111110100" when 4724,
"0001100001110000" when 4725,
"0011110111001101" when 4726,
"0011001011001111" when 4727,
"0000000000001110" when 4728,
"1100110101000011" when 4729,
"1100001000101011" when 4730,
"1110011101110101" when 4731,
"0001111111110011" when 4732,
"0011111101110001" when 4733,
"0010110101001011" when 4734,
"1111011110110101" when 4735,
"1100100010011011" when 4736,
"1100010011011010" when 4737,
"1110111101100010" when 4738,
"0010011011101010" when 4739,
"0011111111111111" when 4740,
"0010011100000001" when 4741,
"1110111101111110" when 4742,
"1100010011100101" when 4743,
"1100100010001100" when 4744,
"1111011110010111" when 4745,
"0010110100110110" when 4746,
"0011111101110101" when 4747,
"0010000000001100" when 4748,
"1110011110010000" when 4749,
"1100001000110011" when 4750,
"1100110100110001" when 4751,
"1111111111110010" when 4752,
"0011001010111101" when 4753,
"0011110111010101" when 4754,
"0001100010001011" when 4755,
"1110000000001101" when 4756,
"1100000010001111" when 4757,
"1101001010110101" when 4758,
"0000100001001011" when 4759,
"0011011101100101" when 4760,
"0011101100100110" when 4761,
"0001000010011110" when 4762,
"1101100100010110" when 4763,
"1100000000000001" when 4764,
"1101100011111111" when 4765,
"0001000010000010" when 4766,
"0011101100011011" when 4767,
"0011011101110100" when 4768,
"0000100001101001" when 4769,
"1101001011001010" when 4770,
"1100000010001011" when 4771,
"1101111111110100" when 4772,
"0001100001110000" when 4773,
"0011110111001101" when 4774,
"0011001011001111" when 4775,
"0000000000001110" when 4776,
"1100110101000011" when 4777,
"1100001000101011" when 4778,
"1110011101110101" when 4779,
"0001111111110011" when 4780,
"0011111101110001" when 4781,
"0010110101001011" when 4782,
"1111011110110101" when 4783,
"1100100010011011" when 4784,
"1100010011011010" when 4785,
"1110111101100010" when 4786,
"0010011011101010" when 4787,
"0011111111111111" when 4788,
"0010011100000001" when 4789,
"1110111101111110" when 4790,
"1100010011100101" when 4791,
"1100100010001100" when 4792,
"1111011110010111" when 4793,
"0010110100110110" when 4794,
"0011111101110101" when 4795,
"0010000000001100" when 4796,
"1110011110010000" when 4797,
"1100001000110011" when 4798,
"1100110100110001" when 4799,
"1111111111110010" when 4800,
"0011001010111101" when 4801,
"0011110111010101" when 4802,
"0001100010001011" when 4803,
"1110000000001101" when 4804,
"1100000010001111" when 4805,
"1101001010110101" when 4806,
"0000100001001011" when 4807,
"0011011101100101" when 4808,
"0011101100100110" when 4809,
"0001000010011111" when 4810,
"1101100100010110" when 4811,
"1100000000000001" when 4812,
"1101100011111111" when 4813,
"0001000010000001" when 4814,
"0011101100011011" when 4815,
"0011011101110100" when 4816,
"0000100001101001" when 4817,
"1101001011001010" when 4818,
"1100000010001011" when 4819,
"1101111111110011" when 4820,
"0001100001101111" when 4821,
"0011110111001101" when 4822,
"0011001011001111" when 4823,
"0000000000001111" when 4824,
"1100110101000011" when 4825,
"1100001000101011" when 4826,
"1110011101110101" when 4827,
"0001111111110010" when 4828,
"0011111101110001" when 4829,
"0010110101001011" when 4830,
"1111011110110101" when 4831,
"1100100010011011" when 4832,
"1100010011011010" when 4833,
"1110111101100001" when 4834,
"0010011011101001" when 4835,
"0011111111111111" when 4836,
"0010011100000001" when 4837,
"1110111101111111" when 4838,
"1100010011100101" when 4839,
"1100100010001100" when 4840,
"1111011110010111" when 4841,
"0010110100110110" when 4842,
"0011111101110101" when 4843,
"0010000000001101" when 4844,
"1110011110010001" when 4845,
"1100001000110011" when 4846,
"1100110100110001" when 4847,
"1111111111110001" when 4848,
"0011001010111101" when 4849,
"0011110111010101" when 4850,
"0001100010001011" when 4851,
"1110000000001110" when 4852,
"1100000010001111" when 4853,
"1101001010110101" when 4854,
"0000100001001011" when 4855,
"0011011101100101" when 4856,
"0011101100100110" when 4857,
"0001000010011111" when 4858,
"1101100100010111" when 4859,
"1100000000000001" when 4860,
"1101100011111111" when 4861,
"0001000010000001" when 4862,
"0011101100011011" when 4863,
"0011011101110100" when 4864,
"0000100001101001" when 4865,
"1101001011001010" when 4866,
"1100000010001011" when 4867,
"1101111111110011" when 4868,
"0001100001101111" when 4869,
"0011110111001101" when 4870,
"0011001011001111" when 4871,
"0000000000001111" when 4872,
"1100110101000011" when 4873,
"1100001000101011" when 4874,
"1110011101110101" when 4875,
"0001111111110010" when 4876,
"0011111101110001" when 4877,
"0010110101001100" when 4878,
"1111011110110101" when 4879,
"1100100010011011" when 4880,
"1100010011011010" when 4881,
"1110111101100001" when 4882,
"0010011011101001" when 4883,
"0011111111111111" when 4884,
"0010011100000010" when 4885,
"1110111101111111" when 4886,
"1100010011100110" when 4887,
"1100100010001100" when 4888,
"1111011110010111" when 4889,
"0010110100110110" when 4890,
"0011111101110101" when 4891,
"0010000000001101" when 4892,
"1110011110010001" when 4893,
"1100001000110011" when 4894,
"1100110100110001" when 4895,
"1111111111110001" when 4896,
"0011001010111100" when 4897,
"0011110111010101" when 4898,
"0001100010001100" when 4899,
"1110000000001110" when 4900,
"1100000010001111" when 4901,
"1101001010110100" when 4902,
"0000100001001011" when 4903,
"0011011101100101" when 4904,
"0011101100100110" when 4905,
"0001000010011111" when 4906,
"1101100100010111" when 4907,
"1100000000000001" when 4908,
"1101100011111110" when 4909,
"0001000010000001" when 4910,
"0011101100011010" when 4911,
"0011011101110100" when 4912,
"0000100001101001" when 4913,
"1101001011001010" when 4914,
"1100000010001011" when 4915,
"1101111111110011" when 4916,
"0001100001101111" when 4917,
"0011110111001101" when 4918,
"0011001011001111" when 4919,
"0000000000001111" when 4920,
"1100110101000100" when 4921,
"1100001000101011" when 4922,
"1110011101110100" when 4923,
"0001111111110010" when 4924,
"0011111101110001" when 4925,
"0010110101001100" when 4926,
"1111011110110101" when 4927,
"1100100010011011" when 4928,
"1100010011011010" when 4929,
"1110111101100001" when 4930,
"0010011011101001" when 4931,
"0011111111111111" when 4932,
"0010011100000010" when 4933,
"1110111101111111" when 4934,
"1100010011100110" when 4935,
"1100100010001100" when 4936,
"1111011110010111" when 4937,
"0010110100110110" when 4938,
"0011111101110101" when 4939,
"0010000000001101" when 4940,
"1110011110010001" when 4941,
"1100001000110011" when 4942,
"1100110100110001" when 4943,
"1111111111110001" when 4944,
"0011001010111100" when 4945,
"0011110111010101" when 4946,
"0001100010001100" when 4947,
"1110000000001110" when 4948,
"1100000010001111" when 4949,
"1101001010110100" when 4950,
"0000100001001011" when 4951,
"0011011101100101" when 4952,
"0011101100100110" when 4953,
"0001000010011111" when 4954,
"1101100100010111" when 4955,
"1100000000000001" when 4956,
"1101100011111110" when 4957,
"0001000010000001" when 4958,
"0011101100011010" when 4959,
"0011011101110100" when 4960,
"0000100001101001" when 4961,
"1101001011001010" when 4962,
"1100000010001011" when 4963,
"1101111111110011" when 4964,
"0001100001101111" when 4965,
"0011110111001101" when 4966,
"0011001011001111" when 4967,
"0000000000001111" when 4968,
"1100110101000100" when 4969,
"1100001000101011" when 4970,
"1110011101110100" when 4971,
"0001111111110010" when 4972,
"0011111101110001" when 4973,
"0010110101001100" when 4974,
"1111011110110101" when 4975,
"1100100010011011" when 4976,
"1100010011011010" when 4977,
"1110111101100001" when 4978,
"0010011011101001" when 4979,
"0011111111111111" when 4980,
"0010011100000010" when 4981,
"1110111101111111" when 4982,
"1100010011100110" when 4983,
"1100100010001100" when 4984,
"1111011110010111" when 4985,
"0010110100110110" when 4986,
"0011111101110101" when 4987,
"0010000000001101" when 4988,
"1110011110010001" when 4989,
"1100001000110011" when 4990,
"1100110100110001" when 4991,
"1111111111110001" when 4992,
"0011001010111100" when 4993,
"0011110111010101" when 4994,
"0001100010001100" when 4995,
"1110000000001110" when 4996,
"1100000010001111" when 4997,
"1101001010110100" when 4998,
"0000100001001011" when 4999,
"0011011101100101" when 5000,
"0011101100100110" when 5001,
"0001000010011111" when 5002,
"1101100100010111" when 5003,
"1100000000000001" when 5004,
"1101100011111110" when 5005,
"0001000010000001" when 5006,
"0011101100011010" when 5007,
"0011011101110100" when 5008,
"0000100001101010" when 5009,
"1101001011001010" when 5010,
"1100000010001011" when 5011,
"1101111111110011" when 5012,
"0001100001101111" when 5013,
"0011110111001101" when 5014,
"0011001011001111" when 5015,
"0000000000001111" when 5016,
"1100110101000100" when 5017,
"1100001000101011" when 5018,
"1110011101110100" when 5019,
"0001111111110010" when 5020,
"0011111101110001" when 5021,
"0010110101001100" when 5022,
"1111011110110110" when 5023,
"1100100010011011" when 5024,
"1100010011011010" when 5025,
"1110111101100001" when 5026,
"0010011011101001" when 5027,
"0011111111111111" when 5028,
"0010011100000010" when 5029,
"1110111101111111" when 5030,
"1100010011100110" when 5031,
"1100100010001100" when 5032,
"1111011110010110" when 5033,
"0010110100110110" when 5034,
"0011111101110101" when 5035,
"0010000000001101" when 5036,
"1110011110010001" when 5037,
"1100001000110011" when 5038,
"1100110100110001" when 5039,
"1111111111110001" when 5040,
"0011001010111100" when 5041,
"0011110111010101" when 5042,
"0001100010001100" when 5043,
"1110000000001110" when 5044,
"1100000010001111" when 5045,
"1101001010110100" when 5046,
"0000100001001010" when 5047,
"0011011101100101" when 5048,
"0011101100100110" when 5049,
"0001000010011111" when 5050,
"1101100100010111" when 5051,
"1100000000000001" when 5052,
"1101100011111110" when 5053,
"0001000010000001" when 5054,
"0011101100011010" when 5055,
"0011011101110100" when 5056,
"0000100001101010" when 5057,
"1101001011001010" when 5058,
"1100000010001011" when 5059,
"1101111111110011" when 5060,
"0001100001101111" when 5061,
"0011110111001101" when 5062,
"0011001011001111" when 5063,
"0000000000001111" when 5064,
"1100110101000100" when 5065,
"1100001000101011" when 5066,
"1110011101110100" when 5067,
"0001111111110010" when 5068,
"0011111101110001" when 5069,
"0010110101001100" when 5070,
"1111011110110110" when 5071,
"1100100010011011" when 5072,
"1100010011011010" when 5073,
"1110111101100001" when 5074,
"0010011011101001" when 5075,
"0011111111111111" when 5076,
"0010011100000010" when 5077,
"1110111101111111" when 5078,
"1100010011100110" when 5079,
"1100100010001100" when 5080,
"1111011110010110" when 5081,
"0010110100110110" when 5082,
"0011111101110101" when 5083,
"0010000000001101" when 5084,
"1110011110010001" when 5085,
"1100001000110011" when 5086,
"1100110100110001" when 5087,
"1111111111110001" when 5088,
"0011001010111100" when 5089,
"0011110111010101" when 5090,
"0001100010001100" when 5091,
"1110000000001110" when 5092,
"1100000010001111" when 5093,
"1101001010110100" when 5094,
"0000100001001010" when 5095,
"0011011101100100" when 5096,
"0011101100100110" when 5097,
"0001000010011111" when 5098,
"1101100100010111" when 5099,
"1100000000000001" when 5100,
"1101100011111110" when 5101,
"0001000010000001" when 5102,
"0011101100011010" when 5103,
"0011011101110100" when 5104,
"0000100001101010" when 5105,
"1101001011001011" when 5106,
"1100000010001011" when 5107,
"1101111111110011" when 5108,
"0001100001101111" when 5109,
"0011110111001101" when 5110,
"0011001011010000" when 5111,
"0000000000001111" when 5112,
"1100110101000100" when 5113,
"1100001000101011" when 5114,
"1110011101110100" when 5115,
"0001111111110010" when 5116,
"0011111101110001" when 5117,
"0010110101001100" when 5118,
"1111011110110110" when 5119,
"1100100010011100" when 5120,
"1100010011011010" when 5121,
"1110111101100001" when 5122,
"0010011011101001" when 5123,
"0011111111111111" when 5124,
"0010011100000010" when 5125,
"1110111101111111" when 5126,
"1100010011100110" when 5127,
"1100100010001100" when 5128,
"1111011110010110" when 5129,
"0010110100110101" when 5130,
"0011111101110101" when 5131,
"0010000000001101" when 5132,
"1110011110010001" when 5133,
"1100001000110011" when 5134,
"1100110100110000" when 5135,
"1111111111110000" when 5136,
"0011001010111100" when 5137,
"0011110111010101" when 5138,
"0001100010001100" when 5139,
"1110000000001110" when 5140,
"1100000010001111" when 5141,
"1101001010110100" when 5142,
"0000100001001010" when 5143,
"0011011101100100" when 5144,
"0011101100100110" when 5145,
"0001000010100000" when 5146,
"1101100100010111" when 5147,
"1100000000000001" when 5148,
"1101100011111110" when 5149,
"0001000010000000" when 5150,
"0011101100011010" when 5151,
"0011011101110100" when 5152,
"0000100001101010" when 5153,
"1101001011001011" when 5154,
"1100000010001011" when 5155,
"1101111111110011" when 5156,
"0001100001101111" when 5157,
"0011110111001101" when 5158,
"0011001011010000" when 5159,
"0000000000010000" when 5160,
"1100110101000100" when 5161,
"1100001000101011" when 5162,
"1110011101110100" when 5163,
"0001111111110010" when 5164,
"0011111101110001" when 5165,
"0010110101001100" when 5166,
"1111011110110110" when 5167,
"1100100010011100" when 5168,
"1100010011011001" when 5169,
"1110111101100000" when 5170,
"0010011011101001" when 5171,
"0011111111111111" when 5172,
"0010011100000010" when 5173,
"1110111110000000" when 5174,
"1100010011100110" when 5175,
"1100100010001011" when 5176,
"1111011110010110" when 5177,
"0010110100110101" when 5178,
"0011111101110101" when 5179,
"0010000000001110" when 5180,
"1110011110010010" when 5181,
"1100001000110011" when 5182,
"1100110100110000" when 5183,
"1111111111110000" when 5184,
"0011001010111100" when 5185,
"0011110111010101" when 5186,
"0001100010001100" when 5187,
"1110000000001111" when 5188,
"1100000010001111" when 5189,
"1101001010110100" when 5190,
"0000100001001010" when 5191,
"0011011101100100" when 5192,
"0011101100100111" when 5193,
"0001000010100000" when 5194,
"1101100100010111" when 5195,
"1100000000000001" when 5196,
"1101100011111110" when 5197,
"0001000010000000" when 5198,
"0011101100011010" when 5199,
"0011011101110101" when 5200,
"0000100001101010" when 5201,
"1101001011001011" when 5202,
"1100000010001011" when 5203,
"1101111111110010" when 5204,
"0001100001101110" when 5205,
"0011110111001101" when 5206,
"0011001011010000" when 5207,
"0000000000010000" when 5208,
"1100110101000100" when 5209,
"1100001000101011" when 5210,
"1110011101110100" when 5211,
"0001111111110001" when 5212,
"0011111101110001" when 5213,
"0010110101001100" when 5214,
"1111011110110110" when 5215,
"1100100010011100" when 5216,
"1100010011011001" when 5217,
"1110111101100000" when 5218,
"0010011011101001" when 5219,
"0011111111111111" when 5220,
"0010011100000010" when 5221,
"1110111110000000" when 5222,
"1100010011100110" when 5223,
"1100100010001011" when 5224,
"1111011110010110" when 5225,
"0010110100110101" when 5226,
"0011111101110101" when 5227,
"0010000000001110" when 5228,
"1110011110010010" when 5229,
"1100001000110011" when 5230,
"1100110100110000" when 5231,
"1111111111110000" when 5232,
"0011001010111100" when 5233,
"0011110111010101" when 5234,
"0001100010001100" when 5235,
"1110000000001111" when 5236,
"1100000010001111" when 5237,
"1101001010110100" when 5238,
"0000100001001010" when 5239,
"0011011101100100" when 5240,
"0011101100100111" when 5241,
"0001000010100000" when 5242,
"1101100100011000" when 5243,
"1100000000000001" when 5244,
"1101100011111110" when 5245,
"0001000010000000" when 5246,
"0011101100011010" when 5247,
"0011011101110101" when 5248,
"0000100001101010" when 5249,
"1101001011001011" when 5250,
"1100000010001011" when 5251,
"1101111111110010" when 5252,
"0001100001101110" when 5253,
"0011110111001101" when 5254,
"0011001011010000" when 5255,
"0000000000010000" when 5256,
"1100110101000100" when 5257,
"1100001000101011" when 5258,
"1110011101110011" when 5259,
"0001111111110001" when 5260,
"0011111101110001" when 5261,
"0010110101001100" when 5262,
"1111011110110110" when 5263,
"1100100010011100" when 5264,
"1100010011011001" when 5265,
"1110111101100000" when 5266,
"0010011011101000" when 5267,
"0011111111111111" when 5268,
"0010011100000010" when 5269,
"1110111110000000" when 5270,
"1100010011100110" when 5271,
"1100100010001011" when 5272,
"1111011110010110" when 5273,
"0010110100110101" when 5274,
"0011111101110101" when 5275,
"0010000000001110" when 5276,
"1110011110010010" when 5277,
"1100001000110011" when 5278,
"1100110100110000" when 5279,
"1111111111110000" when 5280,
"0011001010111100" when 5281,
"0011110111010101" when 5282,
"0001100010001101" when 5283,
"1110000000001111" when 5284,
"1100000010001111" when 5285,
"1101001010110100" when 5286,
"0000100001001010" when 5287,
"0011011101100100" when 5288,
"0011101100100111" when 5289,
"0001000010100000" when 5290,
"1101100100011000" when 5291,
"1100000000000001" when 5292,
"1101100011111101" when 5293,
"0001000010000000" when 5294,
"0011101100011010" when 5295,
"0011011101110101" when 5296,
"0000100001101010" when 5297,
"1101001011001011" when 5298,
"1100000010001011" when 5299,
"1101111111110010" when 5300,
"0001100001101110" when 5301,
"0011110111001101" when 5302,
"0011001011010000" when 5303,
"0000000000010000" when 5304,
"1100110101000100" when 5305,
"1100001000101010" when 5306,
"1110011101110011" when 5307,
"0001111111110001" when 5308,
"0011111101110001" when 5309,
"0010110101001100" when 5310,
"1111011110110110" when 5311,
"1100100010011100" when 5312,
"1100010011011001" when 5313,
"1110111101100000" when 5314,
"0010011011101000" when 5315,
"0011111111111111" when 5316,
"0010011100000011" when 5317,
"1110111110000000" when 5318,
"1100010011100110" when 5319,
"1100100010001011" when 5320,
"1111011110010101" when 5321,
"0010110100110101" when 5322,
"0011111101110101" when 5323,
"0010000000001110" when 5324,
"1110011110010010" when 5325,
"1100001000110011" when 5326,
"1100110100110000" when 5327,
"1111111111110000" when 5328,
"0011001010111100" when 5329,
"0011110111010110" when 5330,
"0001100010001101" when 5331,
"1110000000001111" when 5332,
"1100000010001111" when 5333,
"1101001010110011" when 5334,
"0000100001001010" when 5335,
"0011011101100100" when 5336,
"0011101100100111" when 5337,
"0001000010100000" when 5338,
"1101100100011000" when 5339,
"1100000000000001" when 5340,
"1101100011111101" when 5341,
"0001000010000000" when 5342,
"0011101100011010" when 5343,
"0011011101110101" when 5344,
"0000100001101011" when 5345,
"1101001011001011" when 5346,
"1100000010001010" when 5347,
"1101111111110010" when 5348,
"0001100001101110" when 5349,
"0011110111001101" when 5350,
"0011001011010000" when 5351,
"0000000000010000" when 5352,
"1100110101000100" when 5353,
"1100001000101010" when 5354,
"1110011101110011" when 5355,
"0001111111110001" when 5356,
"0011111101110001" when 5357,
"0010110101001101" when 5358,
"1111011110110111" when 5359,
"1100100010011100" when 5360,
"1100010011011001" when 5361,
"1110111101100000" when 5362,
"0010011011101000" when 5363,
"0011111111111111" when 5364,
"0010011100000011" when 5365,
"1110111110000000" when 5366,
"1100010011100110" when 5367,
"1100100010001011" when 5368,
"1111011110010101" when 5369,
"0010110100110101" when 5370,
"0011111101110110" when 5371,
"0010000000001110" when 5372,
"1110011110010010" when 5373,
"1100001000110011" when 5374,
"1100110100110000" when 5375,
"1111111111110000" when 5376,
"0011001010111100" when 5377,
"0011110111010110" when 5378,
"0001100010001101" when 5379,
"1110000000001111" when 5380,
"1100000010001111" when 5381,
"1101001010110011" when 5382,
"0000100001001001" when 5383,
"0011011101100100" when 5384,
"0011101100100111" when 5385,
"0001000010100000" when 5386,
"1101100100011000" when 5387,
"1100000000000001" when 5388,
"1101100011111101" when 5389,
"0001000010000000" when 5390,
"0011101100011010" when 5391,
"0011011101110101" when 5392,
"0000100001101011" when 5393,
"1101001011001011" when 5394,
"1100000010001010" when 5395,
"1101111111110010" when 5396,
"0001100001101110" when 5397,
"0011110111001101" when 5398,
"0011001011010000" when 5399,
"0000000000010000" when 5400,
"1100110101000100" when 5401,
"1100001000101010" when 5402,
"1110011101110011" when 5403,
"0001111111110001" when 5404,
"0011111101110001" when 5405,
"0010110101001101" when 5406,
"1111011110110111" when 5407,
"1100100010011100" when 5408,
"1100010011011001" when 5409,
"1110111101100000" when 5410,
"0010011011101000" when 5411,
"0011111111111111" when 5412,
"0010011100000011" when 5413,
"1110111110000000" when 5414,
"1100010011100110" when 5415,
"1100100010001011" when 5416,
"1111011110010101" when 5417,
"0010110100110101" when 5418,
"0011111101110110" when 5419,
"0010000000001110" when 5420,
"1110011110010010" when 5421,
"1100001000110011" when 5422,
"1100110100110000" when 5423,
"1111111111110000" when 5424,
"0011001010111011" when 5425,
"0011110111010110" when 5426,
"0001100010001101" when 5427,
"1110000000001111" when 5428,
"1100000010001111" when 5429,
"1101001010110011" when 5430,
"0000100001001001" when 5431,
"0011011101100100" when 5432,
"0011101100100111" when 5433,
"0001000010100000" when 5434,
"1101100100011000" when 5435,
"1100000000000001" when 5436,
"1101100011111101" when 5437,
"0001000010000000" when 5438,
"0011101100011010" when 5439,
"0011011101110101" when 5440,
"0000100001101011" when 5441,
"1101001011001011" when 5442,
"1100000010001010" when 5443,
"1101111111110010" when 5444,
"0001100001101110" when 5445,
"0011110111001101" when 5446,
"0011001011010000" when 5447,
"0000000000010001" when 5448,
"1100110101000101" when 5449,
"1100001000101010" when 5450,
"1110011101110011" when 5451,
"0001111111110001" when 5452,
"0011111101110001" when 5453,
"0010110101001101" when 5454,
"1111011110110111" when 5455,
"1100100010011100" when 5456,
"1100010011011001" when 5457,
"1110111101100000" when 5458,
"0010011011101000" when 5459,
"0011111111111111" when 5460,
"0010011100000011" when 5461,
"1110111110000000" when 5462,
"1100010011100110" when 5463,
"1100100010001011" when 5464,
"1111011110010101" when 5465,
"0010110100110101" when 5466,
"0011111101110110" when 5467,
"0010000000001110" when 5468,
"1110011110010010" when 5469,
"1100001000110011" when 5470,
"1100110100110000" when 5471,
"1111111111101111" when 5472,
"0011001010111011" when 5473,
"0011110111010110" when 5474,
"0001100010001101" when 5475,
"1110000000001111" when 5476,
"1100000010001111" when 5477,
"1101001010110011" when 5478,
"0000100001001001" when 5479,
"0011011101100100" when 5480,
"0011101100100111" when 5481,
"0001000010100001" when 5482,
"1101100100011000" when 5483,
"1100000000000001" when 5484,
"1101100011111101" when 5485,
"0001000001111111" when 5486,
"0011101100011010" when 5487,
"0011011101110101" when 5488,
"0000100001101011" when 5489,
"1101001011001011" when 5490,
"1100000010001010" when 5491,
"1101111111110010" when 5492,
"0001100001101110" when 5493,
"0011110111001101" when 5494,
"0011001011010000" when 5495,
"0000000000010001" when 5496,
"1100110101000101" when 5497,
"1100001000101010" when 5498,
"1110011101110011" when 5499,
"0001111111110001" when 5500,
"0011111101110001" when 5501,
"0010110101001101" when 5502,
"1111011110110111" when 5503,
"1100100010011100" when 5504,
"1100010011011001" when 5505,
"1110111101011111" when 5506,
"0010011011101000" when 5507,
"0011111111111111" when 5508,
"0010011100000011" when 5509,
"1110111110000001" when 5510,
"1100010011100110" when 5511,
"1100100010001011" when 5512,
"1111011110010101" when 5513,
"0010110100110101" when 5514,
"0011111101110110" when 5515,
"0010000000001110" when 5516,
"1110011110010011" when 5517,
"1100001000110011" when 5518,
"1100110100110000" when 5519,
"1111111111101111" when 5520,
"0011001010111011" when 5521,
"0011110111010110" when 5522,
"0001100010001101" when 5523,
"1110000000001111" when 5524,
"1100000010001111" when 5525,
"1101001010110011" when 5526,
"0000100001001001" when 5527,
"0011011101100100" when 5528,
"0011101100100111" when 5529,
"0001000010100001" when 5530,
"1101100100011000" when 5531,
"1100000000000001" when 5532,
"1101100011111101" when 5533,
"0001000001111111" when 5534,
"0011101100011010" when 5535,
"0011011101110101" when 5536,
"0000100001101011" when 5537,
"1101001011001011" when 5538,
"1100000010001010" when 5539,
"1101111111110010" when 5540,
"0001100001101101" when 5541,
"0011110111001101" when 5542,
"0011001011010000" when 5543,
"0000000000010001" when 5544,
"1100110101000101" when 5545,
"1100001000101010" when 5546,
"1110011101110011" when 5547,
"0001111111110000" when 5548,
"0011111101110001" when 5549,
"0010110101001101" when 5550,
"1111011110110111" when 5551,
"1100100010011100" when 5552,
"1100010011011001" when 5553,
"1110111101011111" when 5554,
"0010011011101000" when 5555,
"0011111111111111" when 5556,
"0010011100000011" when 5557,
"1110111110000001" when 5558,
"1100010011100110" when 5559,
"1100100010001011" when 5560,
"1111011110010101" when 5561,
"0010110100110100" when 5562,
"0011111101110110" when 5563,
"0010000000001111" when 5564,
"1110011110010011" when 5565,
"1100001000110011" when 5566,
"1100110100110000" when 5567,
"1111111111101111" when 5568,
"0011001010111011" when 5569,
"0011110111010110" when 5570,
"0001100010001101" when 5571,
"1110000000010000" when 5572,
"1100000010001111" when 5573,
"1101001010110011" when 5574,
"0000100001001001" when 5575,
"0011011101100100" when 5576,
"0011101100100111" when 5577,
"0001000010100001" when 5578,
"1101100100011000" when 5579,
"1100000000000001" when 5580,
"1101100011111101" when 5581,
"0001000001111111" when 5582,
"0011101100011010" when 5583,
"0011011101110101" when 5584,
"0000100001101011" when 5585,
"1101001011001100" when 5586,
"1100000010001010" when 5587,
"1101111111110001" when 5588,
"0001100001101101" when 5589,
"0011110111001101" when 5590,
"0011001011010000" when 5591,
"0000000000010001" when 5592,
"1100110101000101" when 5593,
"1100001000101010" when 5594,
"1110011101110010" when 5595,
"0001111111110000" when 5596,
"0011111101110001" when 5597,
"0010110101001101" when 5598,
"1111011110110111" when 5599,
"1100100010011100" when 5600,
"1100010011011001" when 5601,
"1110111101011111" when 5602,
"0010011011101000" when 5603,
"0011111111111111" when 5604,
"0010011100000011" when 5605,
"1110111110000001" when 5606,
"1100010011100110" when 5607,
"1100100010001011" when 5608,
"1111011110010101" when 5609,
"0010110100110100" when 5610,
"0011111101110110" when 5611,
"0010000000001111" when 5612,
"1110011110010011" when 5613,
"1100001000110011" when 5614,
"1100110100110000" when 5615,
"1111111111101111" when 5616,
"0011001010111011" when 5617,
"0011110111010110" when 5618,
"0001100010001110" when 5619,
"1110000000010000" when 5620,
"1100000010001111" when 5621,
"1101001010110011" when 5622,
"0000100001001001" when 5623,
"0011011101100100" when 5624,
"0011101100100111" when 5625,
"0001000010100001" when 5626,
"1101100100011001" when 5627,
"1100000000000001" when 5628,
"1101100011111101" when 5629,
"0001000001111111" when 5630,
"0011101100011010" when 5631,
"0011011101110101" when 5632,
"0000100001101011" when 5633,
"1101001011001100" when 5634,
"1100000010001010" when 5635,
"1101111111110001" when 5636,
"0001100001101101" when 5637,
"0011110111001101" when 5638,
"0011001011010001" when 5639,
"0000000000010001" when 5640,
"1100110101000101" when 5641,
"1100001000101010" when 5642,
"1110011101110010" when 5643,
"0001111111110000" when 5644,
"0011111101110001" when 5645,
"0010110101001101" when 5646,
"1111011110110111" when 5647,
"1100100010011100" when 5648,
"1100010011011001" when 5649,
"1110111101011111" when 5650,
"0010011011100111" when 5651,
"0011111111111111" when 5652,
"0010011100000011" when 5653,
"1110111110000001" when 5654,
"1100010011100110" when 5655,
"1100100010001011" when 5656,
"1111011110010100" when 5657,
"0010110100110100" when 5658,
"0011111101110110" when 5659,
"0010000000001111" when 5660,
"1110011110010011" when 5661,
"1100001000110011" when 5662,
"1100110100101111" when 5663,
"1111111111101111" when 5664,
"0011001010111011" when 5665,
"0011110111010110" when 5666,
"0001100010001110" when 5667,
"1110000000010000" when 5668,
"1100000010001111" when 5669,
"1101001010110011" when 5670,
"0000100001001000" when 5671,
"0011011101100100" when 5672,
"0011101100100111" when 5673,
"0001000010100001" when 5674,
"1101100100011001" when 5675,
"1100000000000001" when 5676,
"1101100011111100" when 5677,
"0001000001111111" when 5678,
"0011101100011010" when 5679,
"0011011101110101" when 5680,
"0000100001101100" when 5681,
"1101001011001100" when 5682,
"1100000010001010" when 5683,
"1101111111110001" when 5684,
"0001100001101101" when 5685,
"0011110111001101" when 5686,
"0011001011010001" when 5687,
"0000000000010001" when 5688,
"1100110101000101" when 5689,
"1100001000101010" when 5690,
"1110011101110010" when 5691,
"0001111111110000" when 5692,
"0011111101110001" when 5693,
"0010110101001101" when 5694,
"1111011110111000" when 5695,
"1100100010011100" when 5696,
"1100010011011001" when 5697,
"1110111101011111" when 5698,
"0010011011100111" when 5699,
"0011111111111111" when 5700,
"0010011100000100" when 5701,
"1110111110000001" when 5702,
"1100010011100110" when 5703,
"1100100010001011" when 5704,
"1111011110010100" when 5705,
"0010110100110100" when 5706,
"0011111101110110" when 5707,
"0010000000001111" when 5708,
"1110011110010011" when 5709,
"1100001000110011" when 5710,
"1100110100101111" when 5711,
"1111111111101111" when 5712,
"0011001010111011" when 5713,
"0011110111010110" when 5714,
"0001100010001110" when 5715,
"1110000000010000" when 5716,
"1100000010001111" when 5717,
"1101001010110011" when 5718,
"0000100001001000" when 5719,
"0011011101100100" when 5720,
"0011101100100111" when 5721,
"0001000010100001" when 5722,
"1101100100011001" when 5723,
"1100000000000001" when 5724,
"1101100011111100" when 5725,
"0001000001111111" when 5726,
"0011101100011001" when 5727,
"0011011101110101" when 5728,
"0000100001101100" when 5729,
"1101001011001100" when 5730,
"1100000010001010" when 5731,
"1101111111110001" when 5732,
"0001100001101101" when 5733,
"0011110111001101" when 5734,
"0011001011010001" when 5735,
"0000000000010001" when 5736,
"1100110101000101" when 5737,
"1100001000101010" when 5738,
"1110011101110010" when 5739,
"0001111111110000" when 5740,
"0011111101110001" when 5741,
"0010110101001101" when 5742,
"1111011110111000" when 5743,
"1100100010011101" when 5744,
"1100010011011001" when 5745,
"1110111101011111" when 5746,
"0010011011100111" when 5747,
"0011111111111111" when 5748,
"0010011100000100" when 5749,
"1110111110000001" when 5750,
"1100010011100111" when 5751,
"1100100010001011" when 5752,
"1111011110010100" when 5753,
"0010110100110100" when 5754,
"0011111101110110" when 5755,
"0010000000001111" when 5756,
"1110011110010011" when 5757,
"1100001000110011" when 5758,
"1100110100101111" when 5759,
"1111111111101111" when 5760,
"0011001010111011" when 5761,
"0011110111010110" when 5762,
"0001100010001110" when 5763,
"1110000000010000" when 5764,
"1100000010001111" when 5765,
"1101001010110011" when 5766,
"0000100001001000" when 5767,
"0011011101100011" when 5768,
"0011101100100111" when 5769,
"0001000010100001" when 5770,
"1101100100011001" when 5771,
"1100000000000001" when 5772,
"1101100011111100" when 5773,
"0001000001111111" when 5774,
"0011101100011001" when 5775,
"0011011101110101" when 5776,
"0000100001101100" when 5777,
"1101001011001100" when 5778,
"1100000010001010" when 5779,
"1101111111110001" when 5780,
"0001100001101101" when 5781,
"0011110111001101" when 5782,
"0011001011010001" when 5783,
"0000000000010010" when 5784,
"1100110101000101" when 5785,
"1100001000101010" when 5786,
"1110011101110010" when 5787,
"0001111111110000" when 5788,
"0011111101110001" when 5789,
"0010110101001110" when 5790,
"1111011110111000" when 5791,
"1100100010011101" when 5792,
"1100010011011001" when 5793,
"1110111101011111" when 5794,
"0010011011100111" when 5795,
"0011111111111111" when 5796,
"0010011100000100" when 5797,
"1110111110000010" when 5798,
"1100010011100111" when 5799,
"1100100010001010" when 5800,
"1111011110010100" when 5801,
"0010110100110100" when 5802,
"0011111101110110" when 5803,
"0010000000001111" when 5804,
"1110011110010011" when 5805,
"1100001000110011" when 5806,
"1100110100101111" when 5807,
"1111111111101110" when 5808,
"0011001010111011" when 5809,
"0011110111010110" when 5810,
"0001100010001110" when 5811,
"1110000000010000" when 5812,
"1100000010001111" when 5813,
"1101001010110010" when 5814,
"0000100001001000" when 5815,
"0011011101100011" when 5816,
"0011101100100111" when 5817,
"0001000010100010" when 5818,
"1101100100011001" when 5819,
"1100000000000001" when 5820,
"1101100011111100" when 5821,
"0001000001111110" when 5822,
"0011101100011001" when 5823,
"0011011101110110" when 5824,
"0000100001101100" when 5825,
"1101001011001100" when 5826,
"1100000010001010" when 5827,
"1101111111110001" when 5828,
"0001100001101101" when 5829,
"0011110111001101" when 5830,
"0011001011010001" when 5831,
"0000000000010010" when 5832,
"1100110101000101" when 5833,
"1100001000101010" when 5834,
"1110011101110010" when 5835,
"0001111111110000" when 5836,
"0011111101110001" when 5837,
"0010110101001110" when 5838,
"1111011110111000" when 5839,
"1100100010011101" when 5840,
"1100010011011001" when 5841,
"1110111101011110" when 5842,
"0010011011100111" when 5843,
"0011111111111111" when 5844,
"0010011100000100" when 5845,
"1110111110000010" when 5846,
"1100010011100111" when 5847,
"1100100010001010" when 5848,
"1111011110010100" when 5849,
"0010110100110100" when 5850,
"0011111101110110" when 5851,
"0010000000001111" when 5852,
"1110011110010100" when 5853,
"1100001000110100" when 5854,
"1100110100101111" when 5855,
"1111111111101110" when 5856,
"0011001010111011" when 5857,
"0011110111010110" when 5858,
"0001100010001110" when 5859,
"1110000000010000" when 5860,
"1100000010001111" when 5861,
"1101001010110010" when 5862,
"0000100001001000" when 5863,
"0011011101100011" when 5864,
"0011101100100111" when 5865,
"0001000010100010" when 5866,
"1101100100011001" when 5867,
"1100000000000001" when 5868,
"1101100011111100" when 5869,
"0001000001111110" when 5870,
"0011101100011001" when 5871,
"0011011101110110" when 5872,
"0000100001101100" when 5873,
"1101001011001100" when 5874,
"1100000010001010" when 5875,
"1101111111110001" when 5876,
"0001100001101100" when 5877,
"0011110111001100" when 5878,
"0011001011010001" when 5879,
"0000000000010010" when 5880,
"1100110101000101" when 5881,
"1100001000101010" when 5882,
"1110011101110010" when 5883,
"0001111111110000" when 5884,
"0011111101110001" when 5885,
"0010110101001110" when 5886,
"1111011110111000" when 5887,
"1100100010011101" when 5888,
"1100010011011001" when 5889,
"1110111101011110" when 5890,
"0010011011100111" when 5891,
"0011111111111111" when 5892,
"0010011100000100" when 5893,
"1110111110000010" when 5894,
"1100010011100111" when 5895,
"1100100010001010" when 5896,
"1111011110010100" when 5897,
"0010110100110100" when 5898,
"0011111101110110" when 5899,
"0010000000001111" when 5900,
"1110011110010100" when 5901,
"1100001000110100" when 5902,
"1100110100101111" when 5903,
"1111111111101110" when 5904,
"0011001010111011" when 5905,
"0011110111010110" when 5906,
"0001100010001110" when 5907,
"1110000000010000" when 5908,
"1100000010001111" when 5909,
"1101001010110010" when 5910,
"0000100001001000" when 5911,
"0011011101100011" when 5912,
"0011101100100111" when 5913,
"0001000010100010" when 5914,
"1101100100011001" when 5915,
"1100000000000001" when 5916,
"1101100011111100" when 5917,
"0001000001111110" when 5918,
"0011101100011001" when 5919,
"0011011101110110" when 5920,
"0000100001101100" when 5921,
"1101001011001100" when 5922,
"1100000010001010" when 5923,
"1101111111110000" when 5924,
"0001100001101100" when 5925,
"0011110111001100" when 5926,
"0011001011010001" when 5927,
"0000000000010010" when 5928,
"1100110101000101" when 5929,
"1100001000101010" when 5930,
"1110011101110010" when 5931,
"0001111111101111" when 5932,
"0011111101110001" when 5933,
"0010110101001110" when 5934,
"1111011110111000" when 5935,
"1100100010011101" when 5936,
"1100010011011001" when 5937,
"1110111101011110" when 5938,
"0010011011100111" when 5939,
"0011111111111111" when 5940,
"0010011100000100" when 5941,
"1110111110000010" when 5942,
"1100010011100111" when 5943,
"1100100010001010" when 5944,
"1111011110010100" when 5945,
"0010110100110100" when 5946,
"0011111101110110" when 5947,
"0010000000010000" when 5948,
"1110011110010100" when 5949,
"1100001000110100" when 5950,
"1100110100101111" when 5951,
"1111111111101110" when 5952,
"0011001010111010" when 5953,
"0011110111010110" when 5954,
"0001100010001111" when 5955,
"1110000000010001" when 5956,
"1100000010001111" when 5957,
"1101001010110010" when 5958,
"0000100001001000" when 5959,
"0011011101100011" when 5960,
"0011101100100111" when 5961,
"0001000010100010" when 5962,
"1101100100011001" when 5963,
"1100000000000001" when 5964,
"1101100011111100" when 5965,
"0001000001111110" when 5966,
"0011101100011001" when 5967,
"0011011101110110" when 5968,
"0000100001101101" when 5969,
"1101001011001100" when 5970,
"1100000010001010" when 5971,
"1101111111110000" when 5972,
"0001100001101100" when 5973,
"0011110111001100" when 5974,
"0011001011010001" when 5975,
"0000000000010010" when 5976,
"1100110101000110" when 5977,
"1100001000101010" when 5978,
"1110011101110001" when 5979,
"0001111111101111" when 5980,
"0011111101110001" when 5981,
"0010110101001110" when 5982,
"1111011110111000" when 5983,
"1100100010011101" when 5984,
"1100010011011001" when 5985,
"1110111101011110" when 5986,
"0010011011100111" when 5987,
"0011111111111111" when 5988,
"0010011100000100" when 5989,
"1110111110000010" when 5990,
"1100010011100111" when 5991,
"1100100010001010" when 5992,
"1111011110010011" when 5993,
"0010110100110011" when 5994,
"0011111101110110" when 5995,
"0010000000010000" when 5996,
"1110011110010100" when 5997,
"1100001000110100" when 5998,
"1100110100101111" when 5999,
"1111111111101110" when 6000,
"0011001010111010" when 6001,
"0011110111010110" when 6002,
"0001100010001111" when 6003,
"1110000000010001" when 6004,
"1100000010001111" when 6005,
"1101001010110010" when 6006,
"0000100001000111" when 6007,
"0011011101100011" when 6008,
"0011101100101000" when 6009,
"0001000010100010" when 6010,
"1101100100011001" when 6011,
"1100000000000001" when 6012,
"1101100011111100" when 6013,
"0001000001111110" when 6014,
"0011101100011001" when 6015,
"0011011101110110" when 6016,
"0000100001101101" when 6017,
"1101001011001101" when 6018,
"1100000010001010" when 6019,
"1101111111110000" when 6020,
"0001100001101100" when 6021,
"0011110111001100" when 6022,
"0011001011010001" when 6023,
"0000000000010010" when 6024,
"1100110101000110" when 6025,
"1100001000101010" when 6026,
"1110011101110001" when 6027,
"0001111111101111" when 6028,
"0011111101110001" when 6029,
"0010110101001110" when 6030,
"1111011110111001" when 6031,
"1100100010011101" when 6032,
"1100010011011000" when 6033,
"1110111101011110" when 6034,
"0010011011100110" when 6035,
"0011111111111111" when 6036,
"0010011100000100" when 6037,
"1110111110000010" when 6038,
"1100010011100111" when 6039,
"1100100010001010" when 6040,
"1111011110010011" when 6041,
"0010110100110011" when 6042,
"0011111101110110" when 6043,
"0010000000010000" when 6044,
"1110011110010100" when 6045,
"1100001000110100" when 6046,
"1100110100101111" when 6047,
"1111111111101110" when 6048,
"0011001010111010" when 6049,
"0011110111010110" when 6050,
"0001100010001111" when 6051,
"1110000000010001" when 6052,
"1100000010001111" when 6053,
"1101001010110010" when 6054,
"0000100001000111" when 6055,
"0011011101100011" when 6056,
"0011101100101000" when 6057,
"0001000010100010" when 6058,
"1101100100011010" when 6059,
"1100000000000001" when 6060,
"1101100011111100" when 6061,
"0001000001111110" when 6062,
"0011101100011001" when 6063,
"0011011101110110" when 6064,
"0000100001101101" when 6065,
"1101001011001101" when 6066,
"1100000010001010" when 6067,
"1101111111110000" when 6068,
"0001100001101100" when 6069,
"0011110111001100" when 6070,
"0011001011010001" when 6071,
"0000000000010010" when 6072,
"1100110101000110" when 6073,
"1100001000101010" when 6074,
"1110011101110001" when 6075,
"0001111111101111" when 6076,
"0011111101110001" when 6077,
"0010110101001110" when 6078,
"1111011110111001" when 6079,
"1100100010011101" when 6080,
"1100010011011000" when 6081,
"1110111101011110" when 6082,
"0010011011100110" when 6083,
"0011111111111111" when 6084,
"0010011100000101" when 6085,
"1110111110000010" when 6086,
"1100010011100111" when 6087,
"1100100010001010" when 6088,
"1111011110010011" when 6089,
"0010110100110011" when 6090,
"0011111101110110" when 6091,
"0010000000010000" when 6092,
"1110011110010100" when 6093,
"1100001000110100" when 6094,
"1100110100101111" when 6095,
"1111111111101101" when 6096,
"0011001010111010" when 6097,
"0011110111010110" when 6098,
"0001100010001111" when 6099,
"1110000000010001" when 6100,
"1100000010001111" when 6101,
"1101001010110010" when 6102,
"0000100001000111" when 6103,
"0011011101100011" when 6104,
"0011101100101000" when 6105,
"0001000010100010" when 6106,
"1101100100011010" when 6107,
"1100000000000001" when 6108,
"1101100011111011" when 6109,
"0001000001111110" when 6110,
"0011101100011001" when 6111,
"0011011101110110" when 6112,
"0000100001101101" when 6113,
"1101001011001101" when 6114,
"1100000010001010" when 6115,
"1101111111110000" when 6116,
"0001100001101100" when 6117,
"0011110111001100" when 6118,
"0011001011010001" when 6119,
"0000000000010011" when 6120,
"1100110101000110" when 6121,
"1100001000101010" when 6122,
"1110011101110001" when 6123,
"0001111111101111" when 6124,
"0011111101110001" when 6125,
"0010110101001110" when 6126,
"1111011110111001" when 6127,
"1100100010011101" when 6128,
"1100010011011000" when 6129,
"1110111101011110" when 6130,
"0010011011100110" when 6131,
"0011111111111111" when 6132,
"0010011100000101" when 6133,
"1110111110000011" when 6134,
"1100010011100111" when 6135,
"1100100010001010" when 6136,
"1111011110010011" when 6137,
"0010110100110011" when 6138,
"0011111101110110" when 6139,
"0010000000010000" when 6140,
"1110011110010100" when 6141,
"1100001000110100" when 6142,
"1100110100101111" when 6143,
"1111111111101101" when 6144,
"0011001010111010" when 6145,
"0011110111010110" when 6146,
"0001100010001111" when 6147,
"1110000000010001" when 6148,
"1100000010001111" when 6149,
"1101001010110010" when 6150,
"0000100001000111" when 6151,
"0011011101100011" when 6152,
"0011101100101000" when 6153,
"0001000010100011" when 6154,
"1101100100011010" when 6155,
"1100000000000001" when 6156,
"1101100011111011" when 6157,
"0001000001111101" when 6158,
"0011101100011001" when 6159,
"0011011101110110" when 6160,
"0000100001101101" when 6161,
"1101001011001101" when 6162,
"1100000010001010" when 6163,
"1101111111110000" when 6164,
"0001100001101100" when 6165,
"0011110111001100" when 6166,
"0011001011010010" when 6167,
"0000000000010011" when 6168,
"1100110101000110" when 6169,
"1100001000101010" when 6170,
"1110011101110001" when 6171,
"0001111111101111" when 6172,
"0011111101110001" when 6173,
"0010110101001110" when 6174,
"1111011110111001" when 6175,
"1100100010011101" when 6176,
"1100010011011000" when 6177,
"1110111101011101" when 6178,
"0010011011100110" when 6179,
"0011111111111111" when 6180,
"0010011100000101" when 6181,
"1110111110000011" when 6182,
"1100010011100111" when 6183,
"1100100010001010" when 6184,
"1111011110010011" when 6185,
"0010110100110011" when 6186,
"0011111101110110" when 6187,
"0010000000010000" when 6188,
"1110011110010100" when 6189,
"1100001000110100" when 6190,
"1100110100101110" when 6191,
"1111111111101101" when 6192,
"0011001010111010" when 6193,
"0011110111010110" when 6194,
"0001100010001111" when 6195,
"1110000000010001" when 6196,
"1100000010001111" when 6197,
"1101001010110010" when 6198,
"0000100001000111" when 6199,
"0011011101100011" when 6200,
"0011101100101000" when 6201,
"0001000010100011" when 6202,
"1101100100011010" when 6203,
"1100000000000001" when 6204,
"1101100011111011" when 6205,
"0001000001111101" when 6206,
"0011101100011001" when 6207,
"0011011101110110" when 6208,
"0000100001101101" when 6209,
"1101001011001101" when 6210,
"1100000010001010" when 6211,
"1101111111110000" when 6212,
"0001100001101011" when 6213,
"0011110111001100" when 6214,
"0011001011010010" when 6215,
"0000000000010011" when 6216,
"1100110101000110" when 6217,
"1100001000101010" when 6218,
"1110011101110001" when 6219,
"0001111111101111" when 6220,
"0011111101110001" when 6221,
"0010110101001110" when 6222,
"1111011110111001" when 6223,
"1100100010011101" when 6224,
"1100010011011000" when 6225,
"1110111101011101" when 6226,
"0010011011100110" when 6227,
"0011111111111111" when 6228,
"0010011100000101" when 6229,
"1110111110000011" when 6230,
"1100010011100111" when 6231,
"1100100010001010" when 6232,
"1111011110010011" when 6233,
"0010110100110011" when 6234,
"0011111101110110" when 6235,
"0010000000010000" when 6236,
"1110011110010101" when 6237,
"1100001000110100" when 6238,
"1100110100101110" when 6239,
"1111111111101101" when 6240,
"0011001010111010" when 6241,
"0011110111010110" when 6242,
"0001100010001111" when 6243,
"1110000000010001" when 6244,
"1100000010001111" when 6245,
"1101001010110001" when 6246,
"0000100001000111" when 6247,
"0011011101100011" when 6248,
"0011101100101000" when 6249,
"0001000010100011" when 6250,
"1101100100011010" when 6251,
"1100000000000001" when 6252,
"1101100011111011" when 6253,
"0001000001111101" when 6254,
"0011101100011001" when 6255,
"0011011101110110" when 6256,
"0000100001101101" when 6257,
"1101001011001101" when 6258,
"1100000010001010" when 6259,
"1101111111110000" when 6260,
"0001100001101011" when 6261,
"0011110111001100" when 6262,
"0011001011010010" when 6263,
"0000000000010011" when 6264,
"1100110101000110" when 6265,
"1100001000101010" when 6266,
"1110011101110001" when 6267,
"0001111111101111" when 6268,
"0011111101110001" when 6269,
"0010110101001111" when 6270,
"1111011110111001" when 6271,
"1100100010011101" when 6272,
"1100010011011000" when 6273,
"1110111101011101" when 6274,
"0010011011100110" when 6275,
"0011111111111111" when 6276,
"0010011100000101" when 6277,
"1110111110000011" when 6278,
"1100010011100111" when 6279,
"1100100010001010" when 6280,
"1111011110010011" when 6281,
"0010110100110011" when 6282,
"0011111101110110" when 6283,
"0010000000010000" when 6284,
"1110011110010101" when 6285,
"1100001000110100" when 6286,
"1100110100101110" when 6287,
"1111111111101101" when 6288,
"0011001010111010" when 6289,
"0011110111010110" when 6290,
"0001100010010000" when 6291,
"1110000000010010" when 6292,
"1100000010001111" when 6293,
"1101001010110001" when 6294,
"0000100001000111" when 6295,
"0011011101100011" when 6296,
"0011101100101000" when 6297,
"0001000010100011" when 6298,
"1101100100011010" when 6299,
"1100000000000001" when 6300,
"1101100011111011" when 6301,
"0001000001111101" when 6302,
"0011101100011001" when 6303,
"0011011101110110" when 6304,
"0000100001101110" when 6305,
"1101001011001101" when 6306,
"1100000010001010" when 6307,
"1101111111101111" when 6308,
"0001100001101011" when 6309,
"0011110111001100" when 6310,
"0011001011010010" when 6311,
"0000000000010011" when 6312,
"1100110101000110" when 6313,
"1100001000101010" when 6314,
"1110011101110000" when 6315,
"0001111111101110" when 6316,
"0011111101110001" when 6317,
"0010110101001111" when 6318,
"1111011110111010" when 6319,
"1100100010011101" when 6320,
"1100010011011000" when 6321,
"1110111101011101" when 6322,
"0010011011100110" when 6323,
"0011111111111111" when 6324,
"0010011100000101" when 6325,
"1110111110000011" when 6326,
"1100010011100111" when 6327,
"1100100010001010" when 6328,
"1111011110010010" when 6329,
"0010110100110011" when 6330,
"0011111101110110" when 6331,
"0010000000010001" when 6332,
"1110011110010101" when 6333,
"1100001000110100" when 6334,
"1100110100101110" when 6335,
"1111111111101101" when 6336,
"0011001010111010" when 6337,
"0011110111010110" when 6338,
"0001100010010000" when 6339,
"1110000000010010" when 6340,
"1100000010001111" when 6341,
"1101001010110001" when 6342,
"0000100001000110" when 6343,
"0011011101100011" when 6344,
"0011101100101000" when 6345,
"0001000010100011" when 6346,
"1101100100011010" when 6347,
"1100000000000001" when 6348,
"1101100011111011" when 6349,
"0001000001111101" when 6350,
"0011101100011001" when 6351,
"0011011101110110" when 6352,
"0000100001101110" when 6353,
"1101001011001101" when 6354,
"1100000010001010" when 6355,
"1101111111101111" when 6356,
"0001100001101011" when 6357,
"0011110111001100" when 6358,
"0011001011010010" when 6359,
"0000000000010011" when 6360,
"1100110101000110" when 6361,
"1100001000101010" when 6362,
"1110011101110000" when 6363,
"0001111111101110" when 6364,
"0011111101110001" when 6365,
"0010110101001111" when 6366,
"1111011110111010" when 6367,
"1100100010011101" when 6368,
"1100010011011000" when 6369,
"1110111101011101" when 6370,
"0010011011100110" when 6371,
"0011111111111111" when 6372,
"0010011100000101" when 6373,
"1110111110000011" when 6374,
"1100010011100111" when 6375,
"1100100010001010" when 6376,
"1111011110010010" when 6377,
"0010110100110011" when 6378,
"0011111101110110" when 6379,
"0010000000010001" when 6380,
"1110011110010101" when 6381,
"1100001000110100" when 6382,
"1100110100101110" when 6383,
"1111111111101101" when 6384,
"0011001010111010" when 6385,
"0011110111010110" when 6386,
"0001100010010000" when 6387,
"1110000000010010" when 6388,
"1100000010001111" when 6389,
"1101001010110001" when 6390,
"0000100001000110" when 6391,
"0011011101100010" when 6392,
"0011101100101000" when 6393,
"0001000010100011" when 6394,
"1101100100011010" when 6395,
"1100000000000001" when 6396,
"1101100011111011" when 6397,
"0001000001111101" when 6398,
"0011101100011001" when 6399,
"0011011101110110" when 6400,
"0000100001101110" when 6401,
"1101001011001101" when 6402,
"1100000010001010" when 6403,
"1101111111101111" when 6404,
"0001100001101011" when 6405,
"0011110111001100" when 6406,
"0011001011010010" when 6407,
"0000000000010100" when 6408,
"1100110101000110" when 6409,
"1100001000101010" when 6410,
"1110011101110000" when 6411,
"0001111111101110" when 6412,
"0011111101110001" when 6413,
"0010110101001111" when 6414,
"1111011110111010" when 6415,
"1100100010011110" when 6416,
"1100010011011000" when 6417,
"1110111101011101" when 6418,
"0010011011100110" when 6419,
"0011111111111111" when 6420,
"0010011100000101" when 6421,
"1110111110000011" when 6422,
"1100010011100111" when 6423,
"1100100010001010" when 6424,
"1111011110010010" when 6425,
"0010110100110011" when 6426,
"0011111101110110" when 6427,
"0010000000010001" when 6428,
"1110011110010101" when 6429,
"1100001000110100" when 6430,
"1100110100101110" when 6431,
"1111111111101100" when 6432,
"0011001010111010" when 6433,
"0011110111010110" when 6434,
"0001100010010000" when 6435,
"1110000000010010" when 6436,
"1100000010001111" when 6437,
"1101001010110001" when 6438,
"0000100001000110" when 6439,
"0011011101100010" when 6440,
"0011101100101000" when 6441,
"0001000010100011" when 6442,
"1101100100011011" when 6443,
"1100000000000001" when 6444,
"1101100011111011" when 6445,
"0001000001111101" when 6446,
"0011101100011001" when 6447,
"0011011101110111" when 6448,
"0000100001101110" when 6449,
"1101001011001110" when 6450,
"1100000010001010" when 6451,
"1101111111101111" when 6452,
"0001100001101011" when 6453,
"0011110111001100" when 6454,
"0011001011010010" when 6455,
"0000000000010100" when 6456,
"1100110101000110" when 6457,
"1100001000101010" when 6458,
"1110011101110000" when 6459,
"0001111111101110" when 6460,
"0011111101110001" when 6461,
"0010110101001111" when 6462,
"1111011110111010" when 6463,
"1100100010011110" when 6464,
"1100010011011000" when 6465,
"1110111101011101" when 6466,
"0010011011100101" when 6467,
"0011111111111111" when 6468,
"0010011100000101" when 6469,
"1110111110000100" when 6470,
"1100010011100111" when 6471,
"1100100010001001" when 6472,
"1111011110010010" when 6473,
"0010110100110010" when 6474,
"0011111101110110" when 6475,
"0010000000010001" when 6476,
"1110011110010101" when 6477,
"1100001000110100" when 6478,
"1100110100101110" when 6479,
"1111111111101100" when 6480,
"0011001010111001" when 6481,
"0011110111010110" when 6482,
"0001100010010000" when 6483,
"1110000000010010" when 6484,
"1100000010001111" when 6485,
"1101001010110001" when 6486,
"0000100001000110" when 6487,
"0011011101100010" when 6488,
"0011101100101000" when 6489,
"0001000010100100" when 6490,
"1101100100011011" when 6491,
"1100000000000001" when 6492,
"1101100011111010" when 6493,
"0001000001111100" when 6494,
"0011101100011001" when 6495,
"0011011101110111" when 6496,
"0000100001101110" when 6497,
"1101001011001110" when 6498,
"1100000010001010" when 6499,
"1101111111101111" when 6500,
"0001100001101011" when 6501,
"0011110111001100" when 6502,
"0011001011010010" when 6503,
"0000000000010100" when 6504,
"1100110101000111" when 6505,
"1100001000101010" when 6506,
"1110011101110000" when 6507,
"0001111111101110" when 6508,
"0011111101110001" when 6509,
"0010110101001111" when 6510,
"1111011110111010" when 6511,
"1100100010011110" when 6512,
"1100010011011000" when 6513,
"1110111101011100" when 6514,
"0010011011100101" when 6515,
"0011111111111111" when 6516,
"0010011100000110" when 6517,
"1110111110000100" when 6518,
"1100010011100111" when 6519,
"1100100010001001" when 6520,
"1111011110010010" when 6521,
"0010110100110010" when 6522,
"0011111101110110" when 6523,
"0010000000010001" when 6524,
"1110011110010101" when 6525,
"1100001000110100" when 6526,
"1100110100101110" when 6527,
"1111111111101100" when 6528,
"0011001010111001" when 6529,
"0011110111010110" when 6530,
"0001100010010000" when 6531,
"1110000000010010" when 6532,
"1100000010001111" when 6533,
"1101001010110001" when 6534,
"0000100001000110" when 6535,
"0011011101100010" when 6536,
"0011101100101000" when 6537,
"0001000010100100" when 6538,
"1101100100011011" when 6539,
"1100000000000001" when 6540,
"1101100011111010" when 6541,
"0001000001111100" when 6542,
"0011101100011001" when 6543,
"0011011101110111" when 6544,
"0000100001101110" when 6545,
"1101001011001110" when 6546,
"1100000010001010" when 6547,
"1101111111101111" when 6548,
"0001100001101010" when 6549,
"0011110111001100" when 6550,
"0011001011010010" when 6551,
"0000000000010100" when 6552,
"1100110101000111" when 6553,
"1100001000101001" when 6554,
"1110011101110000" when 6555,
"0001111111101110" when 6556,
"0011111101110001" when 6557,
"0010110101001111" when 6558,
"1111011110111010" when 6559,
"1100100010011110" when 6560,
"1100010011011000" when 6561,
"1110111101011100" when 6562,
"0010011011100101" when 6563,
"0011111111111111" when 6564,
"0010011100000110" when 6565,
"1110111110000100" when 6566,
"1100010011101000" when 6567,
"1100100010001001" when 6568,
"1111011110010010" when 6569,
"0010110100110010" when 6570,
"0011111101110110" when 6571,
"0010000000010001" when 6572,
"1110011110010110" when 6573,
"1100001000110100" when 6574,
"1100110100101110" when 6575,
"1111111111101100" when 6576,
"0011001010111001" when 6577,
"0011110111010111" when 6578,
"0001100010010000" when 6579,
"1110000000010010" when 6580,
"1100000010001111" when 6581,
"1101001010110001" when 6582,
"0000100001000110" when 6583,
"0011011101100010" when 6584,
"0011101100101000" when 6585,
"0001000010100100" when 6586,
"1101100100011011" when 6587,
"1100000000000001" when 6588,
"1101100011111010" when 6589,
"0001000001111100" when 6590,
"0011101100011000" when 6591,
"0011011101110111" when 6592,
"0000100001101110" when 6593,
"1101001011001110" when 6594,
"1100000010001010" when 6595,
"1101111111101111" when 6596,
"0001100001101010" when 6597,
"0011110111001100" when 6598,
"0011001011010010" when 6599,
"0000000000010100" when 6600,
"1100110101000111" when 6601,
"1100001000101001" when 6602,
"1110011101110000" when 6603,
"0001111111101110" when 6604,
"0011111101110001" when 6605,
"0010110101001111" when 6606,
"1111011110111010" when 6607,
"1100100010011110" when 6608,
"1100010011011000" when 6609,
"1110111101011100" when 6610,
"0010011011100101" when 6611,
"0011111111111111" when 6612,
"0010011100000110" when 6613,
"1110111110000100" when 6614,
"1100010011101000" when 6615,
"1100100010001001" when 6616,
"1111011110010001" when 6617,
"0010110100110010" when 6618,
"0011111101110110" when 6619,
"0010000000010001" when 6620,
"1110011110010110" when 6621,
"1100001000110100" when 6622,
"1100110100101110" when 6623,
"1111111111101100" when 6624,
"0011001010111001" when 6625,
"0011110111010111" when 6626,
"0001100010010001" when 6627,
"1110000000010010" when 6628,
"1100000010001111" when 6629,
"1101001010110001" when 6630,
"0000100001000110" when 6631,
"0011011101100010" when 6632,
"0011101100101000" when 6633,
"0001000010100100" when 6634,
"1101100100011011" when 6635,
"1100000000000001" when 6636,
"1101100011111010" when 6637,
"0001000001111100" when 6638,
"0011101100011000" when 6639,
"0011011101110111" when 6640,
"0000100001101111" when 6641,
"1101001011001110" when 6642,
"1100000010001010" when 6643,
"1101111111101111" when 6644,
"0001100001101010" when 6645,
"0011110111001100" when 6646,
"0011001011010010" when 6647,
"0000000000010100" when 6648,
"1100110101000111" when 6649,
"1100001000101001" when 6650,
"1110011101101111" when 6651,
"0001111111101110" when 6652,
"0011111101110001" when 6653,
"0010110101001111" when 6654,
"1111011110111011" when 6655,
"1100100010011110" when 6656,
"1100010011011000" when 6657,
"1110111101011100" when 6658,
"0010011011100101" when 6659,
"0011111111111111" when 6660,
"0010011100000110" when 6661,
"1110111110000100" when 6662,
"1100010011101000" when 6663,
"1100100010001001" when 6664,
"1111011110010001" when 6665,
"0010110100110010" when 6666,
"0011111101110110" when 6667,
"0010000000010010" when 6668,
"1110011110010110" when 6669,
"1100001000110100" when 6670,
"1100110100101110" when 6671,
"1111111111101100" when 6672,
"0011001010111001" when 6673,
"0011110111010111" when 6674,
"0001100010010001" when 6675,
"1110000000010011" when 6676,
"1100000010001111" when 6677,
"1101001010110001" when 6678,
"0000100001000101" when 6679,
"0011011101100010" when 6680,
"0011101100101000" when 6681,
"0001000010100100" when 6682,
"1101100100011011" when 6683,
"1100000000000001" when 6684,
"1101100011111010" when 6685,
"0001000001111100" when 6686,
"0011101100011000" when 6687,
"0011011101110111" when 6688,
"0000100001101111" when 6689,
"1101001011001110" when 6690,
"1100000010001010" when 6691,
"1101111111101110" when 6692,
"0001100001101010" when 6693,
"0011110111001100" when 6694,
"0011001011010011" when 6695,
"0000000000010100" when 6696,
"1100110101000111" when 6697,
"1100001000101001" when 6698,
"1110011101101111" when 6699,
"0001111111101101" when 6700,
"0011111101110001" when 6701,
"0010110101010000" when 6702,
"1111011110111011" when 6703,
"1100100010011110" when 6704,
"1100010011011000" when 6705,
"1110111101011100" when 6706,
"0010011011100101" when 6707,
"0011111111111111" when 6708,
"0010011100000110" when 6709,
"1110111110000100" when 6710,
"1100010011101000" when 6711,
"1100100010001001" when 6712,
"1111011110010001" when 6713,
"0010110100110010" when 6714,
"0011111101110110" when 6715,
"0010000000010010" when 6716,
"1110011110010110" when 6717,
"1100001000110100" when 6718,
"1100110100101101" when 6719,
"1111111111101100" when 6720,
"0011001010111001" when 6721,
"0011110111010111" when 6722,
"0001100010010001" when 6723,
"1110000000010011" when 6724,
"1100000010001111" when 6725,
"1101001010110000" when 6726,
"0000100001000101" when 6727,
"0011011101100010" when 6728,
"0011101100101000" when 6729,
"0001000010100100" when 6730,
"1101100100011011" when 6731,
"1100000000000001" when 6732,
"1101100011111010" when 6733,
"0001000001111100" when 6734,
"0011101100011000" when 6735,
"0011011101110111" when 6736,
"0000100001101111" when 6737,
"1101001011001110" when 6738,
"1100000010001010" when 6739,
"1101111111101110" when 6740,
"0001100001101010" when 6741,
"0011110111001100" when 6742,
"0011001011010011" when 6743,
"0000000000010101" when 6744,
"1100110101000111" when 6745,
"1100001000101001" when 6746,
"1110011101101111" when 6747,
"0001111111101101" when 6748,
"0011111101110001" when 6749,
"0010110101010000" when 6750,
"1111011110111011" when 6751,
"1100100010011110" when 6752,
"1100010011011000" when 6753,
"1110111101011100" when 6754,
"0010011011100101" when 6755,
"0011111111111111" when 6756,
"0010011100000110" when 6757,
"1110111110000100" when 6758,
"1100010011101000" when 6759,
"1100100010001001" when 6760,
"1111011110010001" when 6761,
"0010110100110010" when 6762,
"0011111101110110" when 6763,
"0010000000010010" when 6764,
"1110011110010110" when 6765,
"1100001000110100" when 6766,
"1100110100101101" when 6767,
"1111111111101011" when 6768,
"0011001010111001" when 6769,
"0011110111010111" when 6770,
"0001100010010001" when 6771,
"1110000000010011" when 6772,
"1100000010001111" when 6773,
"1101001010110000" when 6774,
"0000100001000101" when 6775,
"0011011101100010" when 6776,
"0011101100101000" when 6777,
"0001000010100100" when 6778,
"1101100100011011" when 6779,
"1100000000000001" when 6780,
"1101100011111010" when 6781,
"0001000001111100" when 6782,
"0011101100011000" when 6783,
"0011011101110111" when 6784,
"0000100001101111" when 6785,
"1101001011001110" when 6786,
"1100000010001010" when 6787,
"1101111111101110" when 6788,
"0001100001101010" when 6789,
"0011110111001100" when 6790,
"0011001011010011" when 6791,
"0000000000010101" when 6792,
"1100110101000111" when 6793,
"1100001000101001" when 6794,
"1110011101101111" when 6795,
"0001111111101101" when 6796,
"0011111101110001" when 6797,
"0010110101010000" when 6798,
"1111011110111011" when 6799,
"1100100010011110" when 6800,
"1100010011011000" when 6801,
"1110111101011011" when 6802,
"0010011011100101" when 6803,
"0011111111111111" when 6804,
"0010011100000110" when 6805,
"1110111110000101" when 6806,
"1100010011101000" when 6807,
"1100100010001001" when 6808,
"1111011110010001" when 6809,
"0010110100110010" when 6810,
"0011111101110110" when 6811,
"0010000000010010" when 6812,
"1110011110010110" when 6813,
"1100001000110100" when 6814,
"1100110100101101" when 6815,
"1111111111101011" when 6816,
"0011001010111001" when 6817,
"0011110111010111" when 6818,
"0001100010010001" when 6819,
"1110000000010011" when 6820,
"1100000010001111" when 6821,
"1101001010110000" when 6822,
"0000100001000101" when 6823,
"0011011101100010" when 6824,
"0011101100101000" when 6825,
"0001000010100101" when 6826,
"1101100100011011" when 6827,
"1100000000000001" when 6828,
"1101100011111010" when 6829,
"0001000001111011" when 6830,
"0011101100011000" when 6831,
"0011011101110111" when 6832,
"0000100001101111" when 6833,
"1101001011001110" when 6834,
"1100000010001010" when 6835,
"1101111111101110" when 6836,
"0001100001101010" when 6837,
"0011110111001100" when 6838,
"0011001011010011" when 6839,
"0000000000010101" when 6840,
"1100110101000111" when 6841,
"1100001000101001" when 6842,
"1110011101101111" when 6843,
"0001111111101101" when 6844,
"0011111101110001" when 6845,
"0010110101010000" when 6846,
"1111011110111011" when 6847,
"1100100010011110" when 6848,
"1100010011010111" when 6849,
"1110111101011011" when 6850,
"0010011011100100" when 6851,
"0011111111111111" when 6852,
"0010011100000110" when 6853,
"1110111110000101" when 6854,
"1100010011101000" when 6855,
"1100100010001001" when 6856,
"1111011110010001" when 6857,
"0010110100110010" when 6858,
"0011111101110110" when 6859,
"0010000000010010" when 6860,
"1110011110010110" when 6861,
"1100001000110100" when 6862,
"1100110100101101" when 6863,
"1111111111101011" when 6864,
"0011001010111001" when 6865,
"0011110111010111" when 6866,
"0001100010010001" when 6867,
"1110000000010011" when 6868,
"1100000010001111" when 6869,
"1101001010110000" when 6870,
"0000100001000101" when 6871,
"0011011101100010" when 6872,
"0011101100101001" when 6873,
"0001000010100101" when 6874,
"1101100100011100" when 6875,
"1100000000000001" when 6876,
"1101100011111010" when 6877,
"0001000001111011" when 6878,
"0011101100011000" when 6879,
"0011011101110111" when 6880,
"0000100001101111" when 6881,
"1101001011001110" when 6882,
"1100000010001010" when 6883,
"1101111111101110" when 6884,
"0001100001101010" when 6885,
"0011110111001100" when 6886,
"0011001011010011" when 6887,
"0000000000010101" when 6888,
"1100110101000111" when 6889,
"1100001000101001" when 6890,
"1110011101101111" when 6891,
"0001111111101101" when 6892,
"0011111101110001" when 6893,
"0010110101010000" when 6894,
"1111011110111011" when 6895,
"1100100010011110" when 6896,
"1100010011010111" when 6897,
"1110111101011011" when 6898,
"0010011011100100" when 6899,
"0011111111111111" when 6900,
"0010011100000111" when 6901,
"1110111110000101" when 6902,
"1100010011101000" when 6903,
"1100100010001001" when 6904,
"1111011110010001" when 6905,
"0010110100110001" when 6906,
"0011111101110110" when 6907,
"0010000000010010" when 6908,
"1110011110010111" when 6909,
"1100001000110100" when 6910,
"1100110100101101" when 6911,
"1111111111101011" when 6912,
"0011001010111001" when 6913,
"0011110111010111" when 6914,
"0001100010010001" when 6915,
"1110000000010011" when 6916,
"1100000010010000" when 6917,
"1101001010110000" when 6918,
"0000100001000101" when 6919,
"0011011101100010" when 6920,
"0011101100101001" when 6921,
"0001000010100101" when 6922,
"1101100100011100" when 6923,
"1100000000000001" when 6924,
"1101100011111001" when 6925,
"0001000001111011" when 6926,
"0011101100011000" when 6927,
"0011011101110111" when 6928,
"0000100001101111" when 6929,
"1101001011001111" when 6930,
"1100000010001010" when 6931,
"1101111111101110" when 6932,
"0001100001101001" when 6933,
"0011110111001100" when 6934,
"0011001011010011" when 6935,
"0000000000010101" when 6936,
"1100110101000111" when 6937,
"1100001000101001" when 6938,
"1110011101101111" when 6939,
"0001111111101101" when 6940,
"0011111101110000" when 6941,
"0010110101010000" when 6942,
"1111011110111011" when 6943,
"1100100010011110" when 6944,
"1100010011010111" when 6945,
"1110111101011011" when 6946,
"0010011011100100" when 6947,
"0011111111111111" when 6948,
"0010011100000111" when 6949,
"1110111110000101" when 6950,
"1100010011101000" when 6951,
"1100100010001001" when 6952,
"1111011110010000" when 6953,
"0010110100110001" when 6954,
"0011111101110110" when 6955,
"0010000000010010" when 6956,
"1110011110010111" when 6957,
"1100001000110100" when 6958,
"1100110100101101" when 6959,
"1111111111101011" when 6960,
"0011001010111001" when 6961,
"0011110111010111" when 6962,
"0001100010010001" when 6963,
"1110000000010011" when 6964,
"1100000010010000" when 6965,
"1101001010110000" when 6966,
"0000100001000100" when 6967,
"0011011101100010" when 6968,
"0011101100101001" when 6969,
"0001000010100101" when 6970,
"1101100100011100" when 6971,
"1100000000000001" when 6972,
"1101100011111001" when 6973,
"0001000001111011" when 6974,
"0011101100011000" when 6975,
"0011011101110111" when 6976,
"0000100001110000" when 6977,
"1101001011001111" when 6978,
"1100000010001010" when 6979,
"1101111111101110" when 6980,
"0001100001101001" when 6981,
"0011110111001100" when 6982,
"0011001011010011" when 6983,
"0000000000010101" when 6984,
"1100110101000111" when 6985,
"1100001000101001" when 6986,
"1110011101101110" when 6987,
"0001111111101101" when 6988,
"0011111101110000" when 6989,
"0010110101010000" when 6990,
"1111011110111100" when 6991,
"1100100010011110" when 6992,
"1100010011010111" when 6993,
"1110111101011011" when 6994,
"0010011011100100" when 6995,
"0011111111111111" when 6996,
"0010011100000111" when 6997,
"1110111110000101" when 6998,
"1100010011101000" when 6999,
"1100100010001001" when 7000,
"1111011110010000" when 7001,
"0010110100110001" when 7002,
"0011111101110110" when 7003,
"0010000000010010" when 7004,
"1110011110010111" when 7005,
"1100001000110100" when 7006,
"1100110100101101" when 7007,
"1111111111101011" when 7008,
"0011001010111000" when 7009,
"0011110111010111" when 7010,
"0001100010010010" when 7011,
"1110000000010011" when 7012,
"1100000010010000" when 7013,
"1101001010110000" when 7014,
"0000100001000100" when 7015,
"0011011101100001" when 7016,
"0011101100101001" when 7017,
"0001000010100101" when 7018,
"1101100100011100" when 7019,
"1100000000000001" when 7020,
"1101100011111001" when 7021,
"0001000001111011" when 7022,
"0011101100011000" when 7023,
"0011011101110111" when 7024,
"0000100001110000" when 7025,
"1101001011001111" when 7026,
"1100000010001010" when 7027,
"1101111111101101" when 7028,
"0001100001101001" when 7029,
"0011110111001100" when 7030,
"0011001011010011" when 7031,
"0000000000010101" when 7032,
"1100110101001000" when 7033,
"1100001000101001" when 7034,
"1110011101101110" when 7035,
"0001111111101100" when 7036,
"0011111101110000" when 7037,
"0010110101010000" when 7038,
"1111011110111100" when 7039,
"1100100010011111" when 7040,
"1100010011010111" when 7041,
"1110111101011011" when 7042,
"0010011011100100" when 7043,
"0011111111111111" when 7044,
"0010011100000111" when 7045,
"1110111110000101" when 7046,
"1100010011101000" when 7047,
"1100100010001001" when 7048,
"1111011110010000" when 7049,
"0010110100110001" when 7050,
"0011111101110110" when 7051,
"0010000000010011" when 7052,
"1110011110010111" when 7053,
"1100001000110100" when 7054,
"1100110100101101" when 7055,
"1111111111101010" when 7056,
"0011001010111000" when 7057,
"0011110111010111" when 7058,
"0001100010010010" when 7059,
"1110000000010100" when 7060,
"1100000010010000" when 7061,
"1101001010110000" when 7062,
"0000100001000100" when 7063,
"0011011101100001" when 7064,
"0011101100101001" when 7065,
"0001000010100101" when 7066,
"1101100100011100" when 7067,
"1100000000000001" when 7068,
"1101100011111001" when 7069,
"0001000001111011" when 7070,
"0011101100011000" when 7071,
"0011011101110111" when 7072,
"0000100001110000" when 7073,
"1101001011001111" when 7074,
"1100000010001010" when 7075,
"1101111111101101" when 7076,
"0001100001101001" when 7077,
"0011110111001011" when 7078,
"0011001011010011" when 7079,
"0000000000010110" when 7080,
"1100110101001000" when 7081,
"1100001000101001" when 7082,
"1110011101101110" when 7083,
"0001111111101100" when 7084,
"0011111101110000" when 7085,
"0010110101010000" when 7086,
"1111011110111100" when 7087,
"1100100010011111" when 7088,
"1100010011010111" when 7089,
"1110111101011011" when 7090,
"0010011011100100" when 7091,
"0011111111111111" when 7092,
"0010011100000111" when 7093,
"1110111110000101" when 7094,
"1100010011101000" when 7095,
"1100100010001000" when 7096,
"1111011110010000" when 7097,
"0010110100110001" when 7098,
"0011111101110110" when 7099,
"0010000000010011" when 7100,
"1110011110010111" when 7101,
"1100001000110101" when 7102,
"1100110100101101" when 7103,
"1111111111101010" when 7104,
"0011001010111000" when 7105,
"0011110111010111" when 7106,
"0001100010010010" when 7107,
"1110000000010100" when 7108,
"1100000010010000" when 7109,
"1101001010110000" when 7110,
"0000100001000100" when 7111,
"0011011101100001" when 7112,
"0011101100101001" when 7113,
"0001000010100101" when 7114,
"1101100100011100" when 7115,
"1100000000000001" when 7116,
"1101100011111001" when 7117,
"0001000001111011" when 7118,
"0011101100011000" when 7119,
"0011011101111000" when 7120,
"0000100001110000" when 7121,
"1101001011001111" when 7122,
"1100000010001010" when 7123,
"1101111111101101" when 7124,
"0001100001101001" when 7125,
"0011110111001011" when 7126,
"0011001011010011" when 7127,
"0000000000010110" when 7128,
"1100110101001000" when 7129,
"1100001000101001" when 7130,
"1110011101101110" when 7131,
"0001111111101100" when 7132,
"0011111101110000" when 7133,
"0010110101010000" when 7134,
"1111011110111100" when 7135,
"1100100010011111" when 7136,
"1100010011010111" when 7137,
"1110111101011010" when 7138,
"0010011011100100" when 7139,
"0011111111111111" when 7140,
"0010011100000111" when 7141,
"1110111110000110" when 7142,
"1100010011101000" when 7143,
"1100100010001000" when 7144,
"1111011110010000" when 7145,
"0010110100110001" when 7146,
"0011111101110110" when 7147,
"0010000000010011" when 7148,
"1110011110010111" when 7149,
"1100001000110101" when 7150,
"1100110100101101" when 7151,
"1111111111101010" when 7152,
"0011001010111000" when 7153,
"0011110111010111" when 7154,
"0001100010010010" when 7155,
"1110000000010100" when 7156,
"1100000010010000" when 7157,
"1101001010101111" when 7158,
"0000100001000100" when 7159,
"0011011101100001" when 7160,
"0011101100101001" when 7161,
"0001000010100110" when 7162,
"1101100100011100" when 7163,
"1100000000000001" when 7164,
"1101100011111001" when 7165,
"0001000001111010" when 7166,
"0011101100011000" when 7167,
"0011011101111000" when 7168,
"0000100001110000" when 7169,
"1101001011001111" when 7170,
"1100000010001010" when 7171,
"1101111111101101" when 7172,
"0001100001101001" when 7173,
"0011110111001011" when 7174,
"0011001011010011" when 7175,
"0000000000010110" when 7176,
"1100110101001000" when 7177,
"1100001000101001" when 7178,
"1110011101101110" when 7179,
"0001111111101100" when 7180,
"0011111101110000" when 7181,
"0010110101010001" when 7182,
"1111011110111100" when 7183,
"1100100010011111" when 7184,
"1100010011010111" when 7185,
"1110111101011010" when 7186,
"0010011011100100" when 7187,
"0011111111111111" when 7188,
"0010011100000111" when 7189,
"1110111110000110" when 7190,
"1100010011101000" when 7191,
"1100100010001000" when 7192,
"1111011110010000" when 7193,
"0010110100110001" when 7194,
"0011111101110110" when 7195,
"0010000000010011" when 7196,
"1110011110010111" when 7197,
"1100001000110101" when 7198,
"1100110100101101" when 7199,
"1111111111101010" when 7200,
"0011001010111000" when 7201,
"0011110111010111" when 7202,
"0001100010010010" when 7203,
"1110000000010100" when 7204,
"1100000010010000" when 7205,
"1101001010101111" when 7206,
"0000100001000100" when 7207,
"0011011101100001" when 7208,
"0011101100101001" when 7209,
"0001000010100110" when 7210,
"1101100100011100" when 7211,
"1100000000000001" when 7212,
"1101100011111001" when 7213,
"0001000001111010" when 7214,
"0011101100011000" when 7215,
"0011011101111000" when 7216,
"0000100001110000" when 7217,
"1101001011001111" when 7218,
"1100000010001010" when 7219,
"1101111111101101" when 7220,
"0001100001101001" when 7221,
"0011110111001011" when 7222,
"0011001011010100" when 7223,
"0000000000010110" when 7224,
"1100110101001000" when 7225,
"1100001000101001" when 7226,
"1110011101101110" when 7227,
"0001111111101100" when 7228,
"0011111101110000" when 7229,
"0010110101010001" when 7230,
"1111011110111100" when 7231,
"1100100010011111" when 7232,
"1100010011010111" when 7233,
"1110111101011010" when 7234,
"0010011011100100" when 7235,
"0011111111111111" when 7236,
"0010011100000111" when 7237,
"1110111110000110" when 7238,
"1100010011101000" when 7239,
"1100100010001000" when 7240,
"1111011110010000" when 7241,
"0010110100110001" when 7242,
"0011111101110110" when 7243,
"0010000000010011" when 7244,
"1110011110011000" when 7245,
"1100001000110101" when 7246,
"1100110100101100" when 7247,
"1111111111101010" when 7248,
"0011001010111000" when 7249,
"0011110111010111" when 7250,
"0001100010010010" when 7251,
"1110000000010100" when 7252,
"1100000010010000" when 7253,
"1101001010101111" when 7254,
"0000100001000100" when 7255,
"0011011101100001" when 7256,
"0011101100101001" when 7257,
"0001000010100110" when 7258,
"1101100100011101" when 7259,
"1100000000000001" when 7260,
"1101100011111001" when 7261,
"0001000001111010" when 7262,
"0011101100011000" when 7263,
"0011011101111000" when 7264,
"0000100001110001" when 7265,
"1101001011001111" when 7266,
"1100000010001010" when 7267,
"1101111111101101" when 7268,
"0001100001101000" when 7269,
"0011110111001011" when 7270,
"0011001011010100" when 7271,
"0000000000010110" when 7272,
"1100110101001000" when 7273,
"1100001000101001" when 7274,
"1110011101101110" when 7275,
"0001111111101100" when 7276,
"0011111101110000" when 7277,
"0010110101010001" when 7278,
"1111011110111101" when 7279,
"1100100010011111" when 7280,
"1100010011010111" when 7281,
"1110111101011010" when 7282,
"0010011011100011" when 7283,
"0011111111111111" when 7284,
"0010011100000111" when 7285,
"1110111110000110" when 7286,
"1100010011101000" when 7287,
"1100100010001000" when 7288,
"1111011110001111" when 7289,
"0010110100110001" when 7290,
"0011111101110110" when 7291,
"0010000000010011" when 7292,
"1110011110011000" when 7293,
"1100001000110101" when 7294,
"1100110100101100" when 7295,
"1111111111101010" when 7296,
"0011001010111000" when 7297,
"0011110111010111" when 7298,
"0001100010010010" when 7299,
"1110000000010100" when 7300,
"1100000010010000" when 7301,
"1101001010101111" when 7302,
"0000100001000011" when 7303,
"0011011101100001" when 7304,
"0011101100101001" when 7305,
"0001000010100110" when 7306,
"1101100100011101" when 7307,
"1100000000000001" when 7308,
"1101100011111000" when 7309,
"0001000001111010" when 7310,
"0011101100011000" when 7311,
"0011011101111000" when 7312,
"0000100001110001" when 7313,
"1101001011001111" when 7314,
"1100000010001010" when 7315,
"1101111111101101" when 7316,
"0001100001101000" when 7317,
"0011110111001011" when 7318,
"0011001011010100" when 7319,
"0000000000010110" when 7320,
"1100110101001000" when 7321,
"1100001000101001" when 7322,
"1110011101101101" when 7323,
"0001111111101100" when 7324,
"0011111101110000" when 7325,
"0010110101010001" when 7326,
"1111011110111101" when 7327,
"1100100010011111" when 7328,
"1100010011010111" when 7329,
"1110111101011010" when 7330,
"0010011011100011" when 7331,
"0011111111111111" when 7332,
"0010011100001000" when 7333,
"1110111110000110" when 7334,
"1100010011101000" when 7335,
"1100100010001000" when 7336,
"1111011110001111" when 7337,
"0010110100110001" when 7338,
"0011111101110110" when 7339,
"0010000000010011" when 7340,
"1110011110011000" when 7341,
"1100001000110101" when 7342,
"1100110100101100" when 7343,
"1111111111101010" when 7344,
"0011001010111000" when 7345,
"0011110111010111" when 7346,
"0001100010010011" when 7347,
"1110000000010100" when 7348,
"1100000010010000" when 7349,
"1101001010101111" when 7350,
"0000100001000011" when 7351,
"0011011101100001" when 7352,
"0011101100101001" when 7353,
"0001000010100110" when 7354,
"1101100100011101" when 7355,
"1100000000000001" when 7356,
"1101100011111000" when 7357,
"0001000001111010" when 7358,
"0011101100011000" when 7359,
"0011011101111000" when 7360,
"0000100001110001" when 7361,
"1101001011010000" when 7362,
"1100000010001010" when 7363,
"1101111111101101" when 7364,
"0001100001101000" when 7365,
"0011110111001011" when 7366,
"0011001011010100" when 7367,
"0000000000010111" when 7368,
"1100110101001000" when 7369,
"1100001000101001" when 7370,
"1110011101101101" when 7371,
"0001111111101100" when 7372,
"0011111101110000" when 7373,
"0010110101010001" when 7374,
"1111011110111101" when 7375,
"1100100010011111" when 7376,
"1100010011010111" when 7377,
"1110111101011010" when 7378,
"0010011011100011" when 7379,
"0011111111111111" when 7380,
"0010011100001000" when 7381,
"1110111110000110" when 7382,
"1100010011101000" when 7383,
"1100100010001000" when 7384,
"1111011110001111" when 7385,
"0010110100110000" when 7386,
"0011111101110110" when 7387,
"0010000000010011" when 7388,
"1110011110011000" when 7389,
"1100001000110101" when 7390,
"1100110100101100" when 7391,
"1111111111101001" when 7392,
"0011001010111000" when 7393,
"0011110111010111" when 7394,
"0001100010010011" when 7395,
"1110000000010101" when 7396,
"1100000010010000" when 7397,
"1101001010101111" when 7398,
"0000100001000011" when 7399,
"0011011101100001" when 7400,
"0011101100101001" when 7401,
"0001000010100110" when 7402,
"1101100100011101" when 7403,
"1100000000000001" when 7404,
"1101100011111000" when 7405,
"0001000001111010" when 7406,
"0011101100010111" when 7407,
"0011011101111000" when 7408,
"0000100001110001" when 7409,
"1101001011010000" when 7410,
"1100000010001010" when 7411,
"1101111111101100" when 7412,
"0001100001101000" when 7413,
"0011110111001011" when 7414,
"0011001011010100" when 7415,
"0000000000010111" when 7416,
"1100110101001000" when 7417,
"1100001000101001" when 7418,
"1110011101101101" when 7419,
"0001111111101011" when 7420,
"0011111101110000" when 7421,
"0010110101010001" when 7422,
"1111011110111101" when 7423,
"1100100010011111" when 7424,
"1100010011010111" when 7425,
"1110111101011010" when 7426,
"0010011011100011" when 7427,
"0011111111111111" when 7428,
"0010011100001000" when 7429,
"1110111110000110" when 7430,
"1100010011101001" when 7431,
"1100100010001000" when 7432,
"1111011110001111" when 7433,
"0010110100110000" when 7434,
"0011111101110110" when 7435,
"0010000000010100" when 7436,
"1110011110011000" when 7437,
"1100001000110101" when 7438,
"1100110100101100" when 7439,
"1111111111101001" when 7440,
"0011001010111000" when 7441,
"0011110111010111" when 7442,
"0001100010010011" when 7443,
"1110000000010101" when 7444,
"1100000010010000" when 7445,
"1101001010101111" when 7446,
"0000100001000011" when 7447,
"0011011101100001" when 7448,
"0011101100101001" when 7449,
"0001000010100110" when 7450,
"1101100100011101" when 7451,
"1100000000000001" when 7452,
"1101100011111000" when 7453,
"0001000001111001" when 7454,
"0011101100010111" when 7455,
"0011011101111000" when 7456,
"0000100001110001" when 7457,
"1101001011010000" when 7458,
"1100000010001010" when 7459,
"1101111111101100" when 7460,
"0001100001101000" when 7461,
"0011110111001011" when 7462,
"0011001011010100" when 7463,
"0000000000010111" when 7464,
"1100110101001000" when 7465,
"1100001000101001" when 7466,
"1110011101101101" when 7467,
"0001111111101011" when 7468,
"0011111101110000" when 7469,
"0010110101010001" when 7470,
"1111011110111101" when 7471,
"1100100010011111" when 7472,
"1100010011010111" when 7473,
"1110111101011001" when 7474,
"0010011011100011" when 7475,
"0011111111111111" when 7476,
"0010011100001000" when 7477,
"1110111110000111" when 7478,
"1100010011101001" when 7479,
"1100100010001000" when 7480,
"1111011110001111" when 7481,
"0010110100110000" when 7482,
"0011111101110110" when 7483,
"0010000000010100" when 7484,
"1110011110011000" when 7485,
"1100001000110101" when 7486,
"1100110100101100" when 7487,
"1111111111101001" when 7488,
"0011001010111000" when 7489,
"0011110111010111" when 7490,
"0001100010010011" when 7491,
"1110000000010101" when 7492,
"1100000010010000" when 7493,
"1101001010101111" when 7494,
"0000100001000011" when 7495,
"0011011101100001" when 7496,
"0011101100101001" when 7497,
"0001000010100111" when 7498,
"1101100100011101" when 7499,
"1100000000000001" when 7500,
"1101100011111000" when 7501,
"0001000001111001" when 7502,
"0011101100010111" when 7503,
"0011011101111000" when 7504,
"0000100001110001" when 7505,
"1101001011010000" when 7506,
"1100000010001010" when 7507,
"1101111111101100" when 7508,
"0001100001101000" when 7509,
"0011110111001011" when 7510,
"0011001011010100" when 7511,
"0000000000010111" when 7512,
"1100110101001000" when 7513,
"1100001000101001" when 7514,
"1110011101101101" when 7515,
"0001111111101011" when 7516,
"0011111101110000" when 7517,
"0010110101010001" when 7518,
"1111011110111101" when 7519,
"1100100010011111" when 7520,
"1100010011010111" when 7521,
"1110111101011001" when 7522,
"0010011011100011" when 7523,
"0011111111111111" when 7524,
"0010011100001000" when 7525,
"1110111110000111" when 7526,
"1100010011101001" when 7527,
"1100100010001000" when 7528,
"1111011110001111" when 7529,
"0010110100110000" when 7530,
"0011111101110110" when 7531,
"0010000000010100" when 7532,
"1110011110011000" when 7533,
"1100001000110101" when 7534,
"1100110100101100" when 7535,
"1111111111101001" when 7536,
"0011001010110111" when 7537,
"0011110111010111" when 7538,
"0001100010010011" when 7539,
"1110000000010101" when 7540,
"1100000010010000" when 7541,
"1101001010101111" when 7542,
"0000100001000011" when 7543,
"0011011101100001" when 7544,
"0011101100101001" when 7545,
"0001000010100111" when 7546,
"1101100100011101" when 7547,
"1100000000000001" when 7548,
"1101100011111000" when 7549,
"0001000001111001" when 7550,
"0011101100010111" when 7551,
"0011011101111000" when 7552,
"0000100001110001" when 7553,
"1101001011010000" when 7554,
"1100000010001010" when 7555,
"1101111111101100" when 7556,
"0001100001101000" when 7557,
"0011110111001011" when 7558,
"0011001011010100" when 7559,
"0000000000010111" when 7560,
"1100110101001001" when 7561,
"1100001000101001" when 7562,
"1110011101101101" when 7563,
"0001111111101011" when 7564,
"0011111101110000" when 7565,
"0010110101010001" when 7566,
"1111011110111101" when 7567,
"1100100010011111" when 7568,
"1100010011010111" when 7569,
"1110111101011001" when 7570,
"0010011011100011" when 7571,
"0011111111111111" when 7572,
"0010011100001000" when 7573,
"1110111110000111" when 7574,
"1100010011101001" when 7575,
"1100100010001000" when 7576,
"1111011110001110" when 7577,
"0010110100110000" when 7578,
"0011111101110110" when 7579,
"0010000000010100" when 7580,
"1110011110011000" when 7581,
"1100001000110101" when 7582,
"1100110100101100" when 7583,
"1111111111101001" when 7584,
"0011001010110111" when 7585,
"0011110111010111" when 7586,
"0001100010010011" when 7587,
"1110000000010101" when 7588,
"1100000010010000" when 7589,
"1101001010101111" when 7590,
"0000100001000011" when 7591,
"0011011101100001" when 7592,
"0011101100101001" when 7593,
"0001000010100111" when 7594,
"1101100100011101" when 7595,
"1100000000000001" when 7596,
"1101100011111000" when 7597,
"0001000001111001" when 7598,
"0011101100010111" when 7599,
"0011011101111000" when 7600,
"0000100001110010" when 7601,
"1101001011010000" when 7602,
"1100000010001010" when 7603,
"1101111111101100" when 7604,
"0001100001100111" when 7605,
"0011110111001011" when 7606,
"0011001011010100" when 7607,
"0000000000010111" when 7608,
"1100110101001001" when 7609,
"1100001000101001" when 7610,
"1110011101101101" when 7611,
"0001111111101011" when 7612,
"0011111101110000" when 7613,
"0010110101010010" when 7614,
"1111011110111110" when 7615,
"1100100010011111" when 7616,
"1100010011010111" when 7617,
"1110111101011001" when 7618,
"0010011011100011" when 7619,
"0011111111111111" when 7620,
"0010011100001000" when 7621,
"1110111110000111" when 7622,
"1100010011101001" when 7623,
"1100100010001000" when 7624,
"1111011110001110" when 7625,
"0010110100110000" when 7626,
"0011111101110110" when 7627,
"0010000000010100" when 7628,
"1110011110011001" when 7629,
"1100001000110101" when 7630,
"1100110100101100" when 7631,
"1111111111101001" when 7632,
"0011001010110111" when 7633,
"0011110111010111" when 7634,
"0001100010010011" when 7635,
"1110000000010101" when 7636,
"1100000010010000" when 7637,
"1101001010101110" when 7638,
"0000100001000010" when 7639,
"0011011101100001" when 7640,
"0011101100101001" when 7641,
"0001000010100111" when 7642,
"1101100100011110" when 7643,
"1100000000000001" when 7644,
"1101100011111000" when 7645,
"0001000001111001" when 7646,
"0011101100010111" when 7647,
"0011011101111000" when 7648,
"0000100001110010" when 7649,
"1101001011010000" when 7650,
"1100000010001010" when 7651,
"1101111111101100" when 7652,
"0001100001100111" when 7653,
"0011110111001011" when 7654,
"0011001011010100" when 7655,
"0000000000010111" when 7656,
"1100110101001001" when 7657,
"1100001000101001" when 7658,
"1110011101101101" when 7659,
"0001111111101011" when 7660,
"0011111101110000" when 7661,
"0010110101010010" when 7662,
"1111011110111110" when 7663,
"1100100010100000" when 7664,
"1100010011010111" when 7665,
"1110111101011001" when 7666,
"0010011011100010" when 7667,
"0011111111111111" when 7668,
"0010011100001000" when 7669,
"1110111110000111" when 7670,
"1100010011101001" when 7671,
"1100100010001000" when 7672,
"1111011110001110" when 7673,
"0010110100110000" when 7674,
"0011111101110110" when 7675,
"0010000000010100" when 7676,
"1110011110011001" when 7677,
"1100001000110101" when 7678,
"1100110100101100" when 7679,
"1111111111101001" when 7680,
"0011001010110111" when 7681,
"0011110111010111" when 7682,
"0001100010010100" when 7683,
"1110000000010101" when 7684,
"1100000010010000" when 7685,
"1101001010101110" when 7686,
"0000100001000010" when 7687,
"0011011101100000" when 7688,
"0011101100101010" when 7689,
"0001000010100111" when 7690,
"1101100100011110" when 7691,
"1100000000000001" when 7692,
"1101100011111000" when 7693,
"0001000001111001" when 7694,
"0011101100010111" when 7695,
"0011011101111000" when 7696,
"0000100001110010" when 7697,
"1101001011010000" when 7698,
"1100000010001010" when 7699,
"1101111111101100" when 7700,
"0001100001100111" when 7701,
"0011110111001011" when 7702,
"0011001011010100" when 7703,
"0000000000011000" when 7704,
"1100110101001001" when 7705,
"1100001000101001" when 7706,
"1110011101101100" when 7707,
"0001111111101011" when 7708,
"0011111101110000" when 7709,
"0010110101010010" when 7710,
"1111011110111110" when 7711,
"1100100010100000" when 7712,
"1100010011010110" when 7713,
"1110111101011001" when 7714,
"0010011011100010" when 7715,
"0011111111111111" when 7716,
"0010011100001001" when 7717,
"1110111110000111" when 7718,
"1100010011101001" when 7719,
"1100100010000111" when 7720,
"1111011110001110" when 7721,
"0010110100110000" when 7722,
"0011111101110110" when 7723,
"0010000000010100" when 7724,
"1110011110011001" when 7725,
"1100001000110101" when 7726,
"1100110100101100" when 7727,
"1111111111101000" when 7728,
"0011001010110111" when 7729,
"0011110111010111" when 7730,
"0001100010010100" when 7731,
"1110000000010101" when 7732,
"1100000010010000" when 7733,
"1101001010101110" when 7734,
"0000100001000010" when 7735,
"0011011101100000" when 7736,
"0011101100101010" when 7737,
"0001000010100111" when 7738,
"1101100100011110" when 7739,
"1100000000000001" when 7740,
"1101100011110111" when 7741,
"0001000001111001" when 7742,
"0011101100010111" when 7743,
"0011011101111001" when 7744,
"0000100001110010" when 7745,
"1101001011010000" when 7746,
"1100000010001010" when 7747,
"1101111111101100" when 7748,
"0001100001100111" when 7749,
"0011110111001011" when 7750,
"0011001011010101" when 7751,
"0000000000011000" when 7752,
"1100110101001001" when 7753,
"1100001000101001" when 7754,
"1110011101101100" when 7755,
"0001111111101011" when 7756,
"0011111101110000" when 7757,
"0010110101010010" when 7758,
"1111011110111110" when 7759,
"1100100010100000" when 7760,
"1100010011010110" when 7761,
"1110111101011001" when 7762,
"0010011011100010" when 7763,
"0011111111111111" when 7764,
"0010011100001001" when 7765,
"1110111110000111" when 7766,
"1100010011101001" when 7767,
"1100100010000111" when 7768,
"1111011110001110" when 7769,
"0010110100110000" when 7770,
"0011111101110110" when 7771,
"0010000000010101" when 7772,
"1110011110011001" when 7773,
"1100001000110101" when 7774,
"1100110100101011" when 7775,
"1111111111101000" when 7776,
"0011001010110111" when 7777,
"0011110111010111" when 7778,
"0001100010010100" when 7779,
"1110000000010110" when 7780,
"1100000010010000" when 7781,
"1101001010101110" when 7782,
"0000100001000010" when 7783,
"0011011101100000" when 7784,
"0011101100101010" when 7785,
"0001000010100111" when 7786,
"1101100100011110" when 7787,
"1100000000000001" when 7788,
"1101100011110111" when 7789,
"0001000001111000" when 7790,
"0011101100010111" when 7791,
"0011011101111001" when 7792,
"0000100001110010" when 7793,
"1101001011010000" when 7794,
"1100000010001010" when 7795,
"1101111111101011" when 7796,
"0001100001100111" when 7797,
"0011110111001011" when 7798,
"0011001011010101" when 7799,
"0000000000011000" when 7800,
"1100110101001001" when 7801,
"1100001000101000" when 7802,
"1110011101101100" when 7803,
"0001111111101010" when 7804,
"0011111101110000" when 7805,
"0010110101010010" when 7806,
"1111011110111110" when 7807,
"1100100010100000" when 7808,
"1100010011010110" when 7809,
"1110111101011000" when 7810,
"0010011011100010" when 7811,
"0011111111111111" when 7812,
"0010011100001001" when 7813,
"1110111110001000" when 7814,
"1100010011101001" when 7815,
"1100100010000111" when 7816,
"1111011110001110" when 7817,
"0010110100101111" when 7818,
"0011111101110111" when 7819,
"0010000000010101" when 7820,
"1110011110011001" when 7821,
"1100001000110101" when 7822,
"1100110100101011" when 7823,
"1111111111101000" when 7824,
"0011001010110111" when 7825,
"0011110111011000" when 7826,
"0001100010010100" when 7827,
"1110000000010110" when 7828,
"1100000010010000" when 7829,
"1101001010101110" when 7830,
"0000100001000010" when 7831,
"0011011101100000" when 7832,
"0011101100101010" when 7833,
"0001000010101000" when 7834,
"1101100100011110" when 7835,
"1100000000000001" when 7836,
"1101100011110111" when 7837,
"0001000001111000" when 7838,
"0011101100010111" when 7839,
"0011011101111001" when 7840,
"0000100001110010" when 7841,
"1101001011010001" when 7842,
"1100000010001001" when 7843,
"1101111111101011" when 7844,
"0001100001100111" when 7845,
"0011110111001011" when 7846,
"0011001011010101" when 7847,
"0000000000011000" when 7848,
"1100110101001001" when 7849,
"1100001000101000" when 7850,
"1110011101101100" when 7851,
"0001111111101010" when 7852,
"0011111101110000" when 7853,
"0010110101010010" when 7854,
"1111011110111110" when 7855,
"1100100010100000" when 7856,
"1100010011010110" when 7857,
"1110111101011000" when 7858,
"0010011011100010" when 7859,
"0011111111111111" when 7860,
"0010011100001001" when 7861,
"1110111110001000" when 7862,
"1100010011101001" when 7863,
"1100100010000111" when 7864,
"1111011110001110" when 7865,
"0010110100101111" when 7866,
"0011111101110111" when 7867,
"0010000000010101" when 7868,
"1110011110011001" when 7869,
"1100001000110101" when 7870,
"1100110100101011" when 7871,
"1111111111101000" when 7872,
"0011001010110111" when 7873,
"0011110111011000" when 7874,
"0001100010010100" when 7875,
"1110000000010110" when 7876,
"1100000010010000" when 7877,
"1101001010101110" when 7878,
"0000100001000010" when 7879,
"0011011101100000" when 7880,
"0011101100101010" when 7881,
"0001000010101000" when 7882,
"1101100100011110" when 7883,
"1100000000000001" when 7884,
"1101100011110111" when 7885,
"0001000001111000" when 7886,
"0011101100010111" when 7887,
"0011011101111001" when 7888,
"0000100001110010" when 7889,
"1101001011010001" when 7890,
"1100000010001001" when 7891,
"1101111111101011" when 7892,
"0001100001100111" when 7893,
"0011110111001011" when 7894,
"0011001011010101" when 7895,
"0000000000011000" when 7896,
"1100110101001001" when 7897,
"1100001000101000" when 7898,
"1110011101101100" when 7899,
"0001111111101010" when 7900,
"0011111101110000" when 7901,
"0010110101010010" when 7902,
"1111011110111110" when 7903,
"1100100010100000" when 7904,
"1100010011010110" when 7905,
"1110111101011000" when 7906,
"0010011011100010" when 7907,
"0011111111111111" when 7908,
"0010011100001001" when 7909,
"1110111110001000" when 7910,
"1100010011101001" when 7911,
"1100100010000111" when 7912,
"1111011110001101" when 7913,
"0010110100101111" when 7914,
"0011111101110111" when 7915,
"0010000000010101" when 7916,
"1110011110011001" when 7917,
"1100001000110101" when 7918,
"1100110100101011" when 7919,
"1111111111101000" when 7920,
"0011001010110111" when 7921,
"0011110111011000" when 7922,
"0001100010010100" when 7923,
"1110000000010110" when 7924,
"1100000010010000" when 7925,
"1101001010101110" when 7926,
"0000100001000001" when 7927,
"0011011101100000" when 7928,
"0011101100101010" when 7929,
"0001000010101000" when 7930,
"1101100100011110" when 7931,
"1100000000000001" when 7932,
"1101100011110111" when 7933,
"0001000001111000" when 7934,
"0011101100010111" when 7935,
"0011011101111001" when 7936,
"0000100001110011" when 7937,
"1101001011010001" when 7938,
"1100000010001001" when 7939,
"1101111111101011" when 7940,
"0001100001100110" when 7941,
"0011110111001011" when 7942,
"0011001011010101" when 7943,
"0000000000011000" when 7944,
"1100110101001001" when 7945,
"1100001000101000" when 7946,
"1110011101101100" when 7947,
"0001111111101010" when 7948,
"0011111101110000" when 7949,
"0010110101010010" when 7950,
"1111011110111111" when 7951,
"1100100010100000" when 7952,
"1100010011010110" when 7953,
"1110111101011000" when 7954,
"0010011011100010" when 7955,
"0011111111111111" when 7956,
"0010011100001001" when 7957,
"1110111110001000" when 7958,
"1100010011101001" when 7959,
"1100100010000111" when 7960,
"1111011110001101" when 7961,
"0010110100101111" when 7962,
"0011111101110111" when 7963,
"0010000000010101" when 7964,
"1110011110011010" when 7965,
"1100001000110101" when 7966,
"1100110100101011" when 7967,
"1111111111101000" when 7968,
"0011001010110111" when 7969,
"0011110111011000" when 7970,
"0001100010010100" when 7971,
"1110000000010110" when 7972,
"1100000010010000" when 7973,
"1101001010101110" when 7974,
"0000100001000001" when 7975,
"0011011101100000" when 7976,
"0011101100101010" when 7977,
"0001000010101000" when 7978,
"1101100100011110" when 7979,
"1100000000000001" when 7980,
"1101100011110111" when 7981,
"0001000001111000" when 7982,
"0011101100010111" when 7983,
"0011011101111001" when 7984,
"0000100001110011" when 7985,
"1101001011010001" when 7986,
"1100000010001001" when 7987,
"1101111111101011" when 7988,
"0001100001100110" when 7989,
"0011110111001011" when 7990,
"0011001011010101" when 7991,
"0000000000011000" when 7992,
"1100110101001001" when 7993,
"1100001000101000" when 7994,
"1110011101101100" when 7995,
"0001111111101010" when 7996,
"0011111101110000" when 7997,
"0010110101010010" when 7998,
"1111011110111111" when 7999,
"1100100010100000" when 8000,
"1100010011010110" when 8001,
"1110111101011000" when 8002,
"0010011011100010" when 8003,
"0011111111111111" when 8004,
"0010011100001001" when 8005,
"1110111110001000" when 8006,
"1100010011101001" when 8007,
"1100100010000111" when 8008,
"1111011110001101" when 8009,
"0010110100101111" when 8010,
"0011111101110111" when 8011,
"0010000000010101" when 8012,
"1110011110011010" when 8013,
"1100001000110101" when 8014,
"1100110100101011" when 8015,
"1111111111100111" when 8016,
"0011001010110111" when 8017,
"0011110111011000" when 8018,
"0001100010010101" when 8019,
"1110000000010110" when 8020,
"1100000010010000" when 8021,
"1101001010101110" when 8022,
"0000100001000001" when 8023,
"0011011101100000" when 8024,
"0011101100101010" when 8025,
"0001000010101000" when 8026,
"1101100100011110" when 8027,
"1100000000000001" when 8028,
"1101100011110111" when 8029,
"0001000001111000" when 8030,
"0011101100010111" when 8031,
"0011011101111001" when 8032,
"0000100001110011" when 8033,
"1101001011010001" when 8034,
"1100000010001001" when 8035,
"1101111111101011" when 8036,
"0001100001100110" when 8037,
"0011110111001011" when 8038,
"0011001011010101" when 8039,
"0000000000011001" when 8040,
"1100110101001010" when 8041,
"1100001000101000" when 8042,
"1110011101101011" when 8043,
"0001111111101010" when 8044,
"0011111101110000" when 8045,
"0010110101010010" when 8046,
"1111011110111111" when 8047,
"1100100010100000" when 8048,
"1100010011010110" when 8049,
"1110111101011000" when 8050,
"0010011011100001" when 8051,
"0011111111111111" when 8052,
"0010011100001001" when 8053,
"1110111110001000" when 8054,
"1100010011101001" when 8055,
"1100100010000111" when 8056,
"1111011110001101" when 8057,
"0010110100101111" when 8058,
"0011111101110111" when 8059,
"0010000000010101" when 8060,
"1110011110011010" when 8061,
"1100001000110101" when 8062,
"1100110100101011" when 8063,
"1111111111100111" when 8064,
"0011001010110110" when 8065,
"0011110111011000" when 8066,
"0001100010010101" when 8067,
"1110000000010110" when 8068,
"1100000010010000" when 8069,
"1101001010101101" when 8070,
"0000100001000001" when 8071,
"0011011101100000" when 8072,
"0011101100101010" when 8073,
"0001000010101000" when 8074,
"1101100100011111" when 8075,
"1100000000000001" when 8076,
"1101100011110111" when 8077,
"0001000001111000" when 8078,
"0011101100010111" when 8079,
"0011011101111001" when 8080,
"0000100001110011" when 8081,
"1101001011010001" when 8082,
"1100000010001001" when 8083,
"1101111111101011" when 8084,
"0001100001100110" when 8085,
"0011110111001011" when 8086,
"0011001011010101" when 8087,
"0000000000011001" when 8088,
"1100110101001010" when 8089,
"1100001000101000" when 8090,
"1110011101101011" when 8091,
"0001111111101010" when 8092,
"0011111101110000" when 8093,
"0010110101010011" when 8094,
"1111011110111111" when 8095,
"1100100010100000" when 8096,
"1100010011010110" when 8097,
"1110111101011000" when 8098,
"0010011011100001" when 8099,
"0011111111111111" when 8100,
"0010011100001010" when 8101,
"1110111110001000" when 8102,
"1100010011101001" when 8103,
"1100100010000111" when 8104,
"1111011110001101" when 8105,
"0010110100101111" when 8106,
"0011111101110111" when 8107,
"0010000000010101" when 8108,
"1110011110011010" when 8109,
"1100001000110101" when 8110,
"1100110100101011" when 8111,
"1111111111100111" when 8112,
"0011001010110110" when 8113,
"0011110111011000" when 8114,
"0001100010010101" when 8115,
"1110000000010110" when 8116,
"1100000010010000" when 8117,
"1101001010101101" when 8118,
"0000100001000001" when 8119,
"0011011101100000" when 8120,
"0011101100101010" when 8121,
"0001000010101000" when 8122,
"1101100100011111" when 8123,
"1100000000000001" when 8124,
"1101100011110110" when 8125,
"0001000001110111" when 8126,
"0011101100010111" when 8127,
"0011011101111001" when 8128,
"0000100001110011" when 8129,
"1101001011010001" when 8130,
"1100000010001001" when 8131,
"1101111111101011" when 8132,
"0001100001100110" when 8133,
"0011110111001011" when 8134,
"0011001011010101" when 8135,
"0000000000011001" when 8136,
"1100110101001010" when 8137,
"1100001000101000" when 8138,
"1110011101101011" when 8139,
"0001111111101001" when 8140,
"0011111101110000" when 8141,
"0010110101010011" when 8142,
"1111011110111111" when 8143,
"1100100010100000" when 8144,
"1100010011010110" when 8145,
"1110111101010111" when 8146,
"0010011011100001" when 8147,
"0011111111111111" when 8148,
"0010011100001010" when 8149,
"1110111110001001" when 8150,
"1100010011101001" when 8151,
"1100100010000111" when 8152,
"1111011110001101" when 8153,
"0010110100101111" when 8154,
"0011111101110111" when 8155,
"0010000000010110" when 8156,
"1110011110011010" when 8157,
"1100001000110101" when 8158,
"1100110100101011" when 8159,
"1111111111100111" when 8160,
"0011001010110110" when 8161,
"0011110111011000" when 8162,
"0001100010010101" when 8163,
"1110000000010111" when 8164,
"1100000010010000" when 8165,
"1101001010101101" when 8166,
"0000100001000001" when 8167,
"0011011101100000" when 8168,
"0011101100101010" when 8169,
"0001000010101001" when 8170,
"1101100100011111" when 8171,
"1100000000000001" when 8172,
"1101100011110110" when 8173,
"0001000001110111" when 8174,
"0011101100010111" when 8175,
"0011011101111001" when 8176,
"0000100001110011" when 8177,
"1101001011010001" when 8178,
"1100000010001001" when 8179,
"1101111111101010" when 8180,
"0001100001100110" when 8181,
"0011110111001011" when 8182,
"0011001011010101" when 8183,
"0000000000011001" when 8184,
"1100110101001010" when 8185,
"1100001000101000" when 8186,
"1110011101101011" when 8187,
"0001111111101001" when 8188,
"0011111101110000" when 8189,
"0010110101010011" when 8190,
"1111011110111111" when 8191,
"0000000000000000" when others;

end Behavioral;